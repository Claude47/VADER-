reg [0:127] wordlist [0:6830] = {"password",
"12345678",
"1q2w3e4r",
"sunshine",
"football",
"computer",
"superman",
"internet",
"iloveyou",
"1qaz2wsx",
"baseball",
"whatever",
"princess",
"abcd1234",
"starwars",
"trustno1",
"jennifer",
"michelle",
"mercedes",
"benjamin",
"11111111",
"samantha",
"victoria",
"asdf1234",
"1234qwer",
"q1w2e3r4",
"elephant",
"garfield",
"jonathan",
"caroline",
"maverick",
"midnight",
"88888888",
"creative",
"cocacola",
"passw0rd",
"blink182",
"danielle",
"scorpion",
"veronica",
"nicholas",
"asdfasdf",
"december",
"patricia",
"security",
"slipknot",
"november",
"jordan23",
"qwertyui",
"carolina",
"hardcore",
"corvette",
"12341234",
"remember",
"qwer1234",
"leonardo",
"snickers",
"williams",
"angelina",
"anderson",
"pakistan",
"marlboro",
"kimberly",
"00000000",
"snowball",
"godzilla",
"hello123",
"champion",
"precious",
"einstein",
"napoleon",
"mountain",
"dolphins",
"fernando",
"87654321",
"paradise",
"motorola",
"bullshit",
"brooklyn",
"qwerty12",
"franklin",
"american",
"platinum",
"icecream",
"darkness",
"cristina",
"colorado",
"steelers",
"serenity",
"mitchell",
"lollipop",
"marshall",
"1qazxsw2",
"12344321",
"startrek",
"business",
"nintendo",
"12qwaszx",
"asdfghjk",
"Password",
"zaq12wsx",
"scotland",
"hercules",
"explorer",
"firebird",
"engineer",
"virginia",
"simpsons",
"angelica",
"isabelle",
"isabella",
"changeme",
"passport",
"infinity",
"courtney",
"scarface",
"pavilion",
"abcdefgh",
"a1b2c3d4",
"harrison",
"spitfire",
"birthday",
"guinness",
"logitech",
"emmanuel",
"11223344",
"goldfish",
"cheyenne",
"testtest",
"stargate",
"anything",
"aaaaaaaa",
"welcome1",
"eternity",
"westside",
"maryjane",
"michael1",
"lawrence",
"kristina",
"kawasaki",
"drowssap",
"blahblah",
"babygirl",
"poohbear",
"florence",
"sapphire",
"hamilton",
"greenday",
"twilight",
"swimming",
"stardust",
"predator",
"penelope",
"michigan",
"margaret",
"brittany",
"shithead",
"redskins",
"pussycat",
"fireball",
"cherokee",
"1234abcd",
"lovelove",
"thailand",
"lasvegas",
"butthead",
"blizzard",
"shamrock",
"bluebird",
"atlantis",
"magnolia",
"juventus",
"diamonds",
"warcraft",
"renegade",
"mohammed",
"shopping",
"savannah",
"giovanni",
"12121212",
"wildcats",
"portugal",
"santiago",
"kathleen",
"clifford",
"55555555",
"rosemary",
"vacation",
"chandler",
"99999999",
"lorraine",
"children",
"beatrice",
"airborne",
"valentin",
"kamikaze",
"software",
"22222222",
"salvador",
"panthers",
"lacrosse",
"charlie1",
"cardinal",
"bluemoon",
"zeppelin",
"rockstar",
"operator",
"dickhead",
"anaconda",
"77777777",
"skittles",
"personal",
"kingkong",
"geronimo",
"robinson",
"kingston",
"hannibal",
"download",
"darkstar",
"sweetpea",
"softball",
"pa55word",
"keyboard",
"darkside",
"assassin",
"vladimir",
"national",
"matthew1",
"brothers",
"warriors",
"universe",
"rush2112",
"mushroom",
"bigdaddy",
"1a2b3c4d",
"ultimate",
"peterpan",
"loverboy",
"truelove",
"trombone",
"madeline",
"gangster",
"dingdong",
"catalina",
"kittycat",
"aquarius",
"patriots",
"ihateyou",
"blessing",
"airplane",
"stingray",
"hellfire",
"guardian",
"flamingo",
"socrates",
"richmond",
"electric",
"thankyou",
"sterling",
"munchkin",
"morpheus",
"imperial",
"goodluck",
"columbia",
"campbell",
"oblivion",
"freedom1",
"valencia",
"spectrum",
"jessica1",
"jeremiah",
"handsome",
"goldberg",
"gabriela",
"anthony1",
"a1234567",
"xxxxxxxx",
"peekaboo",
"montreal",
"kangaroo",
"immortal",
"chocolat",
"thompson",
"research",
"oklahoma",
"mariposa",
"defender",
"applepie",
"squirrel",
"hongkong",
"dinosaur",
"babydoll",
"wolfgang",
"semperfi",
"patience",
"fletcher",
"drpepper",
"creation",
"wordpass",
"passwort",
"original",
"martinez",
"labrador",
"apple123",
"sundance",
"redwings",
"monopoly",
"lionking",
"director",
"44444444",
"sherlock",
"marianne",
"lancelot",
"jeanette",
"cannabis",
"werewolf",
"marathon",
"longhorn",
"happy123",
"brucelee",
"wrangler",
"william1",
"stranger",
"scarlett",
"morrison",
"february",
"fantasia",
"designer",
"bulldogs",
"sullivan",
"saturday",
"pingpong",
"kristine",
"fuckyou1",
"fearless",
"airforce",
"theodore",
"starfish",
"pass1234",
"cinnamon",
"overlord",
"michaela",
"meredith",
"abc12345",
"aardvark",
"Passw0rd",
"trinidad",
"thursday",
"standard",
"pearljam",
"springer",
"ragnarok",
"portland",
"nathalie",
"lemonade",
"lavender",
"gotohell",
"freckles",
"crusader",
"commando",
"clarence",
"cadillac",
"verbatim",
"umbrella",
"splinter",
"register",
"qwert123",
"penguins",
"ncc1701d",
"estrella",
"downtown",
"colombia",
"bollocks",
"69696969",
"showtime",
"qwerasdf",
"mongoose",
"illusion",
"cooldude",
"treasure",
"monalisa",
"justdoit",
"ericsson",
"chelsea1",
"achilles",
"a1s2d3f4",
"veronika",
"test1234",
"sporting",
"papillon",
"juliette",
"fuckyou2",
"firewall",
"cristian",
"cavalier",
"canadian",
"admin123",
"together",
"pa55w0rd",
"halflife",
"formula1",
"thirteen",
"rastaman",
"mustang1",
"cucumber",
"sheridan",
"qqqqqqqq",
"punisher",
"lovelife",
"gretchen",
"chevelle",
"chester1",
"wireless",
"sandiego",
"pokemon1",
"lollypop",
"gorgeous",
"chickens",
"blackman",
"atlantic",
"wildfire",
"waterloo",
"james123",
"homework",
"highland",
"eldorado",
"discover",
"alphabet",
"zaq1xsw2",
"tropical",
"question",
"presario",
"notebook",
"nebraska",
"bullseye",
"valhalla",
"tomorrow",
"richard1",
"positive",
"plymouth",
"patrick1",
"faithful",
"doberman",
"criminal",
"crackers",
"converse",
"casanova",
"attitude",
"66666666",
"scooter1",
"rochelle",
"punkrock",
"kentucky",
"insomnia",
"hooligan",
"gertrude",
"blueeyes",
"terminal",
"poseidon",
"paranoid",
"laurence",
"istanbul",
"frederic",
"doomsday",
"bradford",
"bonehead",
"apollo13",
"westwood",
"satan666",
"reynolds",
"mckenzie",
"magician",
"innocent",
"hotstuff",
"fountain",
"concrete",
"capslock",
"snuggles",
"megadeth",
"medicine",
"jackson1",
"intrepid",
"green123",
"geoffrey",
"dynamite",
"columbus",
"chemical",
"chargers",
"username",
"sherwood",
"moonbeam",
"meowmeow",
"matthias",
"jackson5",
"honolulu",
"diamond1",
"crawford",
"broadway",
"zzzzzzzz",
"whocares",
"svetlana",
"southern",
"pleasure",
"makaveli",
"honeybee",
"francois",
"chicken1",
"bookworm",
"PASSWORD",
"33333333",
"sunlight",
"stallion",
"katerina",
"hedgehog",
"happyday",
"davidson",
"cerberus",
"blackcat",
"arsenal1",
"angel123",
"10101010",
"training",
"republic",
"recovery",
"maradona",
"intruder",
"hermione",
"hastings",
"goldstar",
"fredfred",
"federico",
"deftones",
"blackout",
"1234567a",
"wolfpack",
"thunder1",
"tacobell",
"solution",
"shanghai",
"rootbeer",
"phillips",
"monsters",
"lonewolf",
"keystone",
"johannes",
"grateful",
"continue",
"confused",
"brighton",
"yankees1",
"triangle",
"peterson",
"marianna",
"mandrake",
"inuyasha",
"hardware",
"freebird",
"ferguson",
"dominick",
"bullfrog",
"babylon5",
"13131313",
"zanzibar",
"transfer",
"sparkles",
"shepherd",
"resident",
"property",
"pictures",
"mischief",
"kristian",
"heineken",
"hahahaha",
"eastside",
"daffodil",
"charming",
"billybob",
"adelaide",
"underdog",
"technics",
"samsung1",
"phoenix1",
"musicman",
"marjorie",
"letmein1",
"hospital",
"handball",
"gonzales",
"budapest",
"brandon1",
"alliance",
"adrienne",
"aberdeen",
"thuglife",
"sentinel",
"richards",
"newyork1",
"mortimer",
"marcello",
"magazine",
"infantry",
"hopeless",
"fandango",
"deadhead",
"clarissa",
"christie",
"charlene",
"billyboy",
"bangbang",
"absolute",
"titanium",
"tiger123",
"superior",
"stefanie",
"spaceman",
"somebody",
"sinclair",
"pppppppp",
"mmmmmmmm",
"military",
"loveless",
"karolina",
"fernanda",
"felicity",
"dietcoke",
"brewster",
"babyblue",
"ashleigh",
"14789632",
"whiskers",
"valkyrie",
"superfly",
"strength",
"progress",
"muhammad",
"maryland",
"daughter",
"clarinet",
"chuckles",
"almighty",
"1qaz1qaz",
"sneakers",
"saratoga",
"qawsedrf",
"majestic",
"kingfish",
"japanese",
"graphics",
"flounder",
"coltrane",
"chris123",
"checkers",
"barbados",
"augustus",
"angelika",
"washburn",
"survivor",
"stanford",
"soulmate",
"rasputin",
"pallmall",
"overkill",
"meatloaf",
"lowrider",
"katarina",
"ilovegod",
"heather1",
"hallo123",
"giuseppe",
"eastwood",
"dominion",
"chiquita",
"chipmunk",
"castillo",
"berkeley",
"thinking",
"tarheels",
"seminole",
"pornstar",
"platypus",
"nirvana1",
"mephisto",
"johnjohn",
"gameover",
"fuckface",
"david123",
"darklord",
"cutiepie",
"carnival",
"candyman",
"blowfish",
"ssssssss",
"sandwich",
"sailboat",
"mandarin",
"knuckles",
"jasmine1",
"hardrock",
"boomboom",
"benedict",
"babyface",
"albatros",
"sprinter",
"rolltide",
"r2d2c3po",
"mustangs",
"missouri",
"meridian",
"meatball",
"malaysia",
"killbill",
"illinois",
"gonzalez",
"georgina",
"gargoyle",
"disaster",
"complete",
"claymore",
"chainsaw",
"bluebell",
"98765432",
"wishbone",
"vampires",
"smashing",
"rhiannon",
"rachelle",
"playtime",
"marcella",
"lonestar",
"heritage",
"hayabusa",
"forsaken",
"ferrari1",
"backdoor",
"asshole1",
"11235813",
"yosemite",
"yogibear",
"talisman",
"syracuse",
"randolph",
"raistlin",
"preacher",
"millions",
"metallic",
"madison1",
"dontknow",
"coolcool",
"charisma",
"sinister",
"passpass",
"mohammad",
"mcdonald",
"frontier",
"flipflop",
"eggplant",
"dannyboy",
"daniella",
"chrysler",
"cameron1",
"buckshot",
"arkansas",
"america1",
"12345679",
"romantic",
"robotics",
"redalert",
"megatron",
"mamapapa",
"hyperion",
"gabriel1",
"fuckfuck",
"friendly",
"florida1",
"dreaming",
"doghouse",
"christin",
"brigitte",
"addicted",
"shadow12",
"porkchop",
"negative",
"mistress",
"melissa1",
"jermaine",
"james007",
"francine",
"delphine",
"crystal1",
"chestnut",
"auckland",
"wanderer",
"tomahawk",
"thanatos",
"snoopdog",
"roderick",
"princesa",
"pentagon",
"money123",
"mechanic",
"creature",
"cornwall",
"chadwick",
"calendar",
"abdullah",
"vendetta",
"stephane",
"revolver",
"railroad",
"p4ssw0rd",
"mariners",
"holyshit",
"database",
"bobafett",
"bernardo",
"amethyst",
"advanced",
"whistler",
"slamdunk",
"scrabble",
"roadkill",
"rainbows",
"polopolo",
"obsidian",
"northern",
"learning",
"elements",
"electron",
"customer",
"brisbane",
"baritone",
"amarillo",
"alexandr",
"12301230",
"windmill",
"vanhalen",
"surprise",
"starfire",
"speakers",
"ncc1701e",
"lifetime",
"kittykat",
"fredrick",
"fidelity",
"fabulous",
"everyday",
"coolness",
"concorde",
"catwoman",
"babybaby",
"vodafone",
"traveler",
"rainbow1",
"potatoes",
"pipeline",
"philippe",
"monterey",
"lipstick",
"lakeside",
"insanity",
"fishbone",
"bordeaux",
"21122112",
"windsurf",
"velocity",
"vagabond",
"reloaded",
"raindrop",
"prudence",
"pharmacy",
"peaceful",
"marietta",
"letmein2",
"ladybird",
"internal",
"gigabyte",
"fourteen",
"dolphin1",
"chambers",
"bunghole",
"buckeyes",
"bluefish",
"23232323",
"12369874",
"zerocool",
"wrestler",
"tortoise",
"sysadmin",
"starship",
"qwerty11",
"primrose",
"politics",
"paranoia",
"pancakes",
"overload",
"matthews",
"marriage",
"macaroni",
"jonathon",
"jackjack",
"infinite",
"heinrich",
"graduate",
"goodness",
"godspeed",
"feedback",
"cornelia",
"corleone",
"choochoo",
"chairman",
"butthole",
"buddy123",
"azsxdcfv",
"sleeping",
"pringles",
"power123",
"paradigm",
"nickolas",
"nautilus",
"feathers",
"facebook",
"dragon12",
"brittney",
"aviation",
"19841984",
"10203040",
"wildwood",
"thrasher",
"speedway",
"songbird",
"sickness",
"shannon1",
"screamer",
"monster1",
"mauricio",
"love1234",
"devil666",
"budlight",
"ambrosia",
"adrianna",
"zxcvbnm1",
"windows1",
"toulouse",
"tazmania",
"slapshot",
"ministry",
"mathilde",
"lighting",
"helsinki",
"gateway1",
"fussball",
"frederik",
"flexible",
"festival",
"destiny1",
"daydream",
"coventry",
"constant",
"charles1",
"angeline",
"woodland",
"skinhead",
"sandrine",
"rockford",
"merchant",
"greatest",
"everlast",
"espresso",
"elizabet",
"dddddddd",
"chouchou",
"charlton",
"carlitos",
"blueblue",
"awesome1",
"aspirine",
"12345abc",
"stronger",
"starbuck",
"skeleton",
"scissors",
"reginald",
"redeemer",
"normandy",
"luckydog",
"laserjet",
"just4fun",
"greenbay",
"graffiti",
"doughboy",
"dortmund",
"building",
"bbbbbbbb",
"annabell",
"zimbabwe",
"tunafish",
"thisisit",
"stafford",
"spalding",
"solitude",
"robotech",
"rainbow6",
"qazwsx12",
"pooppoop",
"minister",
"leonidas",
"kirkland",
"integral",
"ilovesex",
"ignatius",
"heavenly",
"gggggggg",
"exchange",
"bulldog1",
"blackdog",
"bearbear",
"winfield",
"westlife",
"thriller",
"spartans",
"sausages",
"printing",
"palmtree",
"opendoor",
"mosquito",
"milkyway",
"laughter",
"klondike",
"kingsley",
"jesus123",
"humphrey",
"hillside",
"hattrick",
"function",
"fighting",
"delaware",
"costello",
"catalyst",
"babylove",
"assholes",
"andersen",
"alexande",
"19891989",
"1234asdf",
"whiplash",
"tiffany1",
"sammy123",
"rockwell",
"reddevil",
"maxwell1",
"gordon24",
"glendale",
"giovanna",
"foxylady",
"fortress",
"favorite",
"doughnut",
"comanche",
"cheshire",
"cherries",
"catarina",
"bertrand",
"barefoot",
"arabella",
"vanguard",
"stephen1",
"rhapsody",
"reckless",
"pumpkin1",
"powerful",
"painting",
"nocturne",
"nickname",
"mynameis",
"mikemike",
"llllllll",
"leighton",
"kkkkkkkk",
"johnston",
"holidays",
"handyman",
"fuckoff1",
"front242",
"flamenco",
"escalade",
"division",
"covenant",
"cannibal",
"annmarie",
"alcatraz",
"11112222",
"wwwwwwww",
"wildcard",
"whitesox",
"vincent1",
"thornton",
"survival",
"sprocket",
"somerset",
"skorpion",
"services",
"restless",
"pumpkins",
"meathead",
"lucky123",
"licorice",
"language",
"jackass1",
"infiniti",
"gamecube",
"flanders",
"disciple",
"diplomat",
"crescent",
"catholic",
"capoeira",
"browning",
"biscuits",
"alexalex",
"P@ssw0rd",
"Jennifer",
"19861986",
"winston1",
"violator",
"super123",
"straight",
"sorcerer",
"sidekick",
"shredder",
"schubert",
"prestige",
"peter123",
"nonsense",
"mulligan",
"moneyman",
"matchbox",
"marauder",
"longhair",
"lisalisa",
"kayleigh",
"islander",
"genesis1",
"gardenia",
"gabriele",
"edmonton",
"downhill",
"digital1",
"cromwell",
"chowchow",
"carebear",
"vanessa1",
"terrapin",
"stockton",
"smoothie",
"seahawks",
"rebecca1",
"rangers1",
"puppydog",
"marigold",
"gregorio",
"gangbang",
"dutchess",
"daylight",
"clueless",
"calamity",
"beefcake",
"aquarium",
"anathema",
"ambition",
"19821982",
"wildlife",
"snowbird",
"qwerqwer",
"prospect",
"natalie1",
"lockdown",
"italiano",
"irishman",
"infamous",
"hydrogen",
"hartford",
"goodyear",
"generals",
"garrison",
"foxhound",
"entrance",
"eighteen",
"diamante",
"daedalus",
"cocktail",
"caligula",
"borabora",
"behemoth",
"balloons",
"bachelor",
"waterman",
"teenager",
"spanking",
"soccer10",
"sergeant",
"seashell",
"seahorse",
"riffraff",
"possible",
"pinnacle",
"nostromo",
"latitude",
"kevin123",
"invasion",
"hibiscus",
"hallmark",
"envision",
"charcoal",
"blue1234",
"antelope",
"aircraft",
"123456aa",
"viktoria",
"stripper",
"stefania",
"smirnoff",
"seraphim",
"ronaldo7",
"reporter",
"raiders1",
"nineteen",
"monolith",
"memories",
"memorial",
"massacre",
"honduras",
"goofball",
"fullmoon",
"forever1",
"elefante",
"doorknob",
"dipstick",
"commerce",
"carousel",
"callisto",
"berenice",
"asdfzxcv",
"alex1234",
"Welcome1",
"19871987",
"wormwood",
"starstar",
"sexygirl",
"rosewood",
"roadster",
"rapunzel",
"prisoner",
"prescott",
"pizza123",
"phillies",
"phantom1",
"perfect1",
"pasadena",
"optimist",
"master12",
"junkmail",
"inspiron",
"hhhhhhhh",
"griffith",
"golfball",
"forester",
"euphoria",
"england1",
"death666",
"conquest",
"clitoris",
"cartoons",
"buckaroo",
"bluejays",
"violence",
"testpass",
"terrence",
"temporal",
"teamwork",
"spencer1",
"shipping",
"roosters",
"prophecy",
"popcorn1",
"playmate",
"panorama",
"p0o9i8u7",
"landmark",
"johnson1",
"iverson3",
"instinct",
"infected",
"honeydew",
"document",
"deadline",
"cowboys1",
"climbing",
"bubbles1",
"bluestar",
"bathroom",
"anamaria",
"25802580",
"24682468",
"whiteboy",
"titleist",
"tiberius",
"retarded",
"palomino",
"outsider",
"oooooooo",
"musician",
"michelin",
"hyacinth",
"gatorade",
"fuzzball",
"everyone",
"delirium",
"daisy123",
"critical",
"cordelia",
"capitals",
"caliente",
"bobdylan",
"Michelle",
"1a2s3d4f",
"19781978",
"voltaire",
"thedoors",
"special1",
"southpaw",
"soccer12",
"ruthless",
"reaction",
"qazwsxed",
"portable",
"passcode",
"official",
"mindless",
"masamune",
"lalalala",
"holloway",
"hairball",
"dirtbike",
"dilligaf",
"clippers",
"chicago1",
"caldwell",
"agent007",
"19831983",
"19801980",
"19751975",
"warrior1",
"vertical",
"timeless",
"thegreat",
"spelling",
"slippery",
"rrrrrrrr",
"ricochet",
"protocol",
"producer",
"penguin1",
"p455w0rd",
"olivetti",
"oliveira",
"metalica",
"mannheim",
"mandingo",
"magellan",
"machines",
"lovebird",
"jason123",
"inflames",
"headache",
"godbless",
"gemstone",
"ffffffff",
"cyclones",
"colonial",
"claudius",
"bulgaria",
"brunette",
"bradshaw",
"bastards",
"basement",
"acapulco",
"25252525",
"12312312",
"zachary1",
"yingyang",
"workshop",
"trueblue",
"sycamore",
"stigmata",
"sabrina1",
"riccardo",
"playboy1",
"override",
"music123",
"mortgage",
"meandyou",
"macdaddy",
"knockers",
"kisskiss",
"jjjjjjjj",
"hysteria",
"forgiven",
"distance",
"cosworth",
"coconuts",
"carlisle",
"asdfjkl;",
"31415926",
"21212121",
"yokohama",
"tommy123",
"sheepdog",
"seinfeld",
"sabotage",
"pressure",
"pinetree",
"pavement",
"oriental",
"offshore",
"netscape",
"michaels",
"mash4077",
"mallorca",
"junkyard",
"johncena",
"jakejake",
"hawthorn",
"hawaiian",
"frenchie",
"fishing1",
"fastball",
"deathrow",
"calimero",
"breakout",
"black123",
"bismarck",
"alkaline",
"zxcv1234",
"tryagain",
"thatcher",
"stampede",
"scheisse",
"sayonara",
"passions",
"nothing1",
"nameless",
"mysterio",
"monkey12",
"millwall",
"megabyte",
"mccarthy",
"magister",
"madhouse",
"liverpoo",
"laetitia",
"jennings",
"holstein",
"freefall",
"flawless",
"ebenezer",
"divinity",
"delpiero",
"chastity",
"charlott",
"carlotta",
"buchanan",
"bradley1",
"aventura",
"asdffdsa",
"19741974",
"zildjian",
"wargames",
"vvvvvvvv",
"unicorns",
"tenerife",
"tasmania",
"symphony",
"splendid",
"sonyvaio",
"snapshot",
"saunders",
"sarajevo",
"reverend",
"polaroid",
"perfecto",
"nokia123",
"natasha1",
"mystical",
"melanie1",
"material",
"maddison",
"landlord",
"juvenile",
"goodwill",
"goldwing",
"gilberto",
"gandalf1",
"fuckthis",
"flapjack",
"flamengo",
"finnegan",
"fabienne",
"erection",
"clemente",
"caterina",
"capetown",
"antonio1",
"angelito",
"accounts",
"abstract",
"19911991",
"19761976",
"01234567",
"vincenzo",
"townsend",
"soccer11",
"smithers",
"shooting",
"shitshit",
"senators",
"redbaron",
"percival",
"painless",
"myfamily",
"mongolia",
"miroslav",
"macarena",
"lakewood",
"killer12",
"incoming",
"immanuel",
"hometown",
"homeless",
"giordano",
"genocide",
"enforcer",
"dispatch",
"codename",
"cccccccc",
"caramelo",
"callaway",
"calculus",
"brian123",
"blessed1",
"attorney",
"asteroid",
"academia",
"12131415",
"yamahar1",
"tricolor",
"terrance",
"summer99",
"stirling",
"stamford",
"stairway",
"soldiers",
"shitface",
"scorpio1",
"principe",
"pizzahut",
"patricio",
"passwerd",
"mulberry",
"luscious",
"lifeline",
"legoland",
"kickflip",
"kennwort",
"kathrine",
"josefina",
"jesus777",
"hellsing",
"drummond",
"delldell",
"cupcakes",
"claudine",
"ciaociao",
"christia",
"cashmere",
"carthage",
"bookmark",
"bartlett",
"alphonse",
"Benjamin",
"51505150",
"woodside",
"vaseline",
"trinity1",
"toxicity",
"tommyboy",
"ticktock",
"teachers",
"strategy",
"stephens",
"snowdrop",
"smeghead",
"shutdown",
"sexysexy",
"popsicle",
"petersen",
"oscar123",
"maryanne",
"magicman",
"kingking",
"identity",
"icehouse",
"hannover",
"glorious",
"forgetit",
"fishtank",
"epiphone",
"elevator",
"elegance",
"drumline",
"devilman",
"delivery",
"chrissie",
"carnaval",
"caffeine",
"bukowski",
"brownies",
"bearcats",
"akatsuki",
"19941994",
"woofwoof",
"virginie",
"untitled",
"tttttttt",
"timothy1",
"stickman",
"starlite",
"smarties",
"oxymoron",
"oleander",
"ncc1701a",
"muhammed",
"morphine",
"mobydick",
"meltdown",
"medieval",
"mahogany",
"magic123",
"longshot",
"lockheed",
"livewire",
"lakeland",
"kenworth",
"interpol",
"hunter12",
"hibernia",
"helpdesk",
"godofwar",
"fishhead",
"ethernet",
"duracell",
"crystals",
"colossus",
"besiktas",
"backlash",
"academic",
"abnormal",
"19901990",
"violetta",
"vineyard",
"terrible",
"suburban",
"stocking",
"snuffles",
"sideways",
"schwartz",
"salasana",
"rosalind",
"purchase",
"practice",
"poiuytre",
"piramide",
"montrose",
"molly123",
"maximus1",
"mammamia",
"lunchbox",
"lonesome",
"limerick",
"liberty1",
"ignition",
"homebrew",
"harry123",
"greenman",
"godsmack",
"firefire",
"daniel12",
"cricket1",
"contract",
"conflict",
"comeback",
"coldplay",
"believer",
"beaumont",
"angelita",
"23456789",
"woodward",
"wolverin",
"wellness",
"swingers",
"solstice",
"scratchy",
"rockport",
"redlight",
"puppy123",
"paulette",
"panther1",
"overtime",
"nazareth",
"mudvayne",
"movement",
"miracles",
"mike1234",
"maserati",
"marbella",
"kiwikiwi",
"jurassic",
"infernal",
"hereford",
"goodtime",
"goodlife",
"goodgirl",
"gamecock",
"gabriell",
"friends1",
"ferreira",
"ethiopia",
"dionysus",
"deadpool",
"christos",
"chauncey",
"castaway",
"carefree",
"burnside",
"borussia",
"bohemian",
"blackice",
"bigmouth",
"baptiste",
"augustin",
"asdfg123",
"alistair",
"advocate",
"adgjmptw",
"acoustic",
"Princess",
"19811981",
"11221122",
"youandme",
"vinicius",
"vauxhall",
"tyler123",
"terminus",
"surround",
"soccer13",
"sexylady",
"sessions",
"scirocco",
"schiller",
"schedule",
"rosebud1",
"regional",
"radiance",
"pioneers",
"phantasy",
"peaches1",
"p@ssw0rd",
"neutrino",
"kendrick",
"hogwarts",
"heinlein",
"guitarra",
"gillette",
"germania",
"flowers1",
"fighters",
"fastback",
"fabrizio",
"exercise",
"envelope",
"element1",
"eeeeeeee",
"doraemon",
"diabetes",
"damascus",
"coronado",
"cashflow",
"cardigan",
"blackboy",
"bitchass",
"backpack",
"anakonda",
"Victoria",
"911turbo",
"19851985",
"19721972",
"water123",
"viscount",
"violette",
"undertow",
"teacher1",
"success1",
"stephani",
"redstone",
"premiere",
"planning",
"paramore",
"packers1",
"nitrogen",
"natascha",
"moonwalk",
"maurizio",
"marzipan",
"mandolin",
"mamamama",
"maintain",
"macgyver",
"ludacris",
"loredana",
"killkill",
"justice1",
"jailbird",
"goodnews",
"freshman",
"firestar",
"eleonora",
"dragon11",
"domenico",
"discreet",
"crossbow",
"choppers",
"betrayed",
"bernhard",
"basilisk",
"antigone",
"alterego",
"alhambra",
"aerobics",
"Superman",
"20012001",
"1million",
"yyyyyyyy",
"woodruff",
"vampire1",
"tequiero",
"sunnyboy",
"specialk",
"sorrento",
"reliance",
"q2w3e4r5",
"proverbs",
"playgirl",
"pentium4",
"pedigree",
"partners",
"orange12",
"observer",
"nnnnnnnn",
"newworld",
"moriarty",
"minotaur",
"location",
"knockout",
"knickers",
"jeffrey1",
"hellyeah",
"greentea",
"goodgood",
"germany1",
"gasoline",
"flashman",
"fatality",
"emiliano",
"ellipsis",
"disorder",
"deadlock",
"davidoff",
"couscous",
"congress",
"cleaning",
"clarkson",
"charlie2",
"ceramics",
"casandra",
"cambodia",
"bigmoney",
"backbone",
"74108520",
"24681012",
"24242424",
"19881988",
"whatwhat",
"watching",
"tomatoes",
"tiramisu",
"tiberian",
"thurston",
"spinning",
"slippers",
"simon123",
"response",
"reindeer",
"porsche1",
"panchito",
"montana1",
"mayfield",
"marquise",
"manifest",
"magnetic",
"lovelace",
"lesbians",
"joystick",
"industry",
"gulliver",
"ganymede",
"galactic",
"esoteric",
"dropdead",
"drinking",
"devildog",
"copeland",
"christop",
"cheerios",
"chatting",
"changeit",
"cerulean",
"cabernet",
"bionicle",
"baltazar",
"amoremio",
"alpha123",
"alleycat",
"accident",
"19771977",
"123mudar",
"tingting",
"thething",
"testing1",
"tallulah",
"symmetry",
"summer69",
"smartass",
"shadow11",
"salesman",
"rushmore",
"resource",
"pregnant",
"pleasant",
"plankton",
"pendulum",
"paterson",
"partizan",
"olympics",
"networks",
"mystique",
"mckinley",
"mcgregor",
"maxpower",
"livelife",
"kokakola",
"katherin",
"julianna",
"jeannine",
"horseman",
"homeland",
"holiday1",
"hennessy",
"guesswho",
"greywolf",
"gilligan",
"gallardo",
"freewill",
"francis1",
"fordf150",
"fantomas",
"dutchman",
"drummer1",
"dementia",
"berliner",
"20002000",
"19951995",
"woodwork",
"winifred",
"welcome2",
"waterboy",
"troopers",
"theodora",
"sometime",
"russell1",
"roadking",
"rifleman",
"raymond1",
"qwerty13",
"priyanka",
"private1",
"pizzaman",
"phantasm",
"pathetic",
"nicotine",
"mollydog",
"minstrel",
"matthieu",
"maria123",
"lebron23",
"lakers24",
"kitty123",
"kindness",
"hatfield",
"getmoney",
"general1",
"forsythe",
"fontaine",
"feelgood",
"evidence",
"erickson",
"enter123",
"downfall",
"deadwood",
"crazyman",
"citation",
"calliope",
"broccoli",
"bleeding",
"bergkamp",
"asmodeus",
"artistic",
"antilles",
"anteater",
"anhyeuem",
"aaaa1111",
"Sunshine",
"Jonathan",
"19731973",
"19691969",
"wrinkles",
"trumpet1",
"triplets",
"sunnyday",
"summer12",
"students",
"start123",
"sopranos",
"siberian",
"shetland",
"sheppard",
"scrapper",
"schooner",
"pershing",
"parasite",
"pantera1",
"palmetto",
"overture",
"odysseus",
"noisette",
"narayana",
"nakamura",
"mediator",
"mcintosh",
"mazda626",
"marykate",
"manpower",
"malamute",
"justin12",
"jeronimo",
"jeremias",
"jamaican",
"imperium",
"humberto",
"hotmail1",
"hoosiers",
"goldmine",
"futurama",
"elisabet",
"dumpling",
"dragster",
"dragon13",
"dominica",
"dominate",
"dictator",
"cookbook",
"concerto",
"christel",
"beholder",
"babushka",
"autobahn",
"anywhere",
"acidburn",
"abhishek",
"z1x2c3v4",
"whiteout",
"topolino",
"thousand",
"thorsten",
"symantec",
"stanley1",
"splatter",
"sonysony",
"schaefer",
"reddwarf",
"position",
"popopopo",
"pikapika",
"piercing",
"pasquale",
"neighbor",
"mireille",
"lovesick",
"loverman",
"london12",
"lockwood",
"kowalski",
"kerberos",
"kellyann",
"jimmy123",
"jayhawks",
"innuendo",
"ilovemom",
"iiiiiiii",
"houston1",
"horrible",
"himalaya",
"highlife",
"hetfield",
"graphite",
"funnyman",
"f00tball",
"epiphany",
"elvis123",
"discount",
"danny123",
"consumer",
"chouette",
"chinchin",
"chinaman",
"calderon",
"bullhead",
"brussels",
"brasilia",
"bobby123",
"bellevue",
"bagpipes",
"aurelius",
"altitude",
"aloysius",
"alabama1",
"affinity",
"abcdefg1",
"20102010",
"09876543",
"zxasqw12",
"winnipeg",
"ultraman",
"treefrog",
"tigercat",
"taratara",
"tactical",
"system32",
"swastika",
"skipper1",
"searcher",
"reserved",
"redbeard",
"realtime",
"pyramids",
"provider",
"projects",
"poontang",
"pinecone",
"pericles",
"paradiso",
"parabola",
"overflow",
"mazdarx7",
"marybeth",
"marriott",
"madalena",
"loophole",
"lonsdale",
"lingerie",
"libertad",
"lavalamp",
"joselito",
"joker123",
"jerrylee",
"jamboree",
"interest",
"imissyou",
"hugoboss",
"holahola",
"heythere",
"hehehehe",
"hangover",
"guerrero",
"greatone",
"gianluca",
"gardener",
"gangsta1",
"exorcist",
"dressage",
"dominic1",
"dodgeram",
"cummings",
"christen",
"callahan",
"calcutta",
"burberry",
"betrayal",
"atkinson",
"athletic",
"arachnid",
"amaranth",
"algernon",
"alastair",
"absinthe",
"01020304",
"zoomzoom",
"watchman",
"vanilla1",
"trouble1",
"tortilla",
"squadron",
"smile123",
"skylight",
"ricardo1",
"reliable",
"recorder",
"provence",
"porsche9",
"piedmont",
"patches1",
"overdose",
"nightman",
"mymother",
"monument",
"medicina",
"madonna1",
"longtime",
"lolololo",
"lokiloki",
"laughing",
"kerrigan",
"jeopardy",
"ibelieve",
"houghton",
"horsemen",
"hologram",
"hideaway",
"hawaii50",
"handicap",
"hamsters",
"georgia1",
"freddie1",
"forklift",
"finished",
"dorothea",
"devotion",
"conchita",
"classics",
"chopper1",
"buffalo1",
"bubba123",
"bigballs",
"barnyard",
"baphomet",
"badlands",
"asterisk",
"arcangel",
"20022002",
"19971997",
"whoknows",
"trousers",
"tranquil",
"toriamos",
"temppass",
"teardrop",
"superboy",
"srinivas",
"snowman1",
"shortcut",
"shocking",
"senha123",
"scranton",
"sandoval",
"roseanne",
"red12345",
"prospero",
"products",
"papamama",
"outdoors",
"nemesis1",
"nagasaki",
"mousepad",
"modeling",
"microlab",
"makeitso",
"lalakers",
"kakaroto",
"investor",
"insecure",
"humanoid",
"holiness",
"helpless",
"germaine",
"freefree",
"francais",
"firebolt",
"filipino",
"federica",
"falstaff",
"eleven11",
"dominant",
"diabolic",
"deadbeat",
"crockett",
"crazycat",
"composer",
"coleslaw",
"cascades",
"bretagne",
"breaking",
"bluenose",
"bisexual",
"billions",
"billbill",
"beckham7",
"avengers",
"assembly",
"asasasas",
"allstars",
"alakazam",
"activate",
"Pa55word",
"Computer",
"zerozero",
"vigilant",
"verygood",
"truffles",
"tigerman",
"thankgod",
"telefono",
"summoner",
"suicidal",
"strummer",
"stiletto",
"squeaker",
"sithlord",
"showcase",
"serenade",
"rotation",
"rockhard",
"quintana",
"pacifica",
"omsairam",
"newhouse",
"nacional",
"muenchen",
"morrigan",
"michael2",
"memememe",
"maximize",
"marino13",
"marciano",
"loveable",
"lakeview",
"kenneth1",
"ilikepie",
"historia",
"hiawatha",
"freeport",
"flathead",
"faulkner",
"endymion",
"emirates",
"dreamers",
"dragon69",
"district",
"dietrich",
"clemence",
"claudia1",
"cellular",
"catherin",
"carmella",
"burgundy",
"brother1",
"blooming",
"bigboobs",
"beachbum",
"barbara1",
"backyard",
"backward",
"babybear",
"argonaut",
"appleton",
"aguilera",
"Nicholas",
"Michael1",
"1qazzaq1",
"13243546",
"12qw34er",
"123456ab",
"zaragoza",
"woodcock",
"wisteria",
"westlake",
"victoire",
"trapdoor",
"tigereye",
"thetruth",
"testicle",
"student1",
"sprinkle",
"silencer",
"scottish",
"richelle",
"religion",
"queenbee",
"physical",
"pedersen",
"paperboy",
"nikolaus",
"murderer",
"montague",
"milagros",
"mercutio",
"mercurio",
"mcknight",
"maxpayne",
"manager1",
"mamacita",
"lucretia",
"lol12345",
"laura123",
"kusanagi",
"katmandu",
"julianne",
"joseluis",
"jiujitsu",
"jeanpaul",
"infrared",
"humanity",
"honeypot",
"honeybun",
"herkules",
"hawkeyes",
"gregory1",
"geometry",
"friedman",
"freiheit",
"firework",
"elbereth",
"dragon99",
"dollface",
"devilish",
"democrat",
"darkmoon",
"crackpot",
"costanza",
"consuelo",
"clarisse",
"citibank",
"cingular",
"chrystal",
"channing",
"carvalho",
"brownie1",
"bluebear",
"billyjoe",
"benedikt",
"beaufort",
"batman12",
"barnabas",
"baracuda",
"armitage",
"alcapone",
"adrianne",
"a1a2a3a4",
"Internet",
"Football",
"yourself",
"yorktown",
"yeahyeah",
"valdemar",
"unlocked",
"twinkles",
"trujillo",
"torrents",
"tonyhawk",
"tanzania",
"takedown",
"takamine",
"stitches",
"standing",
"srilanka",
"sparhawk",
"slowpoke",
"shoelace",
"service1",
"senorita",
"seashore",
"roulette",
"rocky123",
"radiator",
"problems",
"platform",
"parallax",
"nepenthe",
"moonmoon",
"lovehate",
"komputer",
"intrigue",
"interact",
"galloway",
"fullback",
"fuckhead",
"fairview",
"divorced",
"disabled",
"defiance",
"deeznutz",
"daniel01",
"cookies1",
"cheating",
"boarding",
"baseline",
"baldrick",
"apollo11",
"aluminum",
"19931993",
"19791979",
"woodwind",
"woodbury",
"watchdog",
"vikings1",
"tribunal",
"toreador",
"thinkpad",
"thebeach",
"terrific",
"teaching",
"stringer",
"souvenir",
"sombrero",
"sk8board",
"shuriken",
"shotokan",
"shinichi",
"scooters",
"regiment",
"rainfall",
"qwerty78",
"pistache",
"pianoman",
"overseas",
"orthodox",
"monorail",
"minemine",
"milhouse",
"mermaids",
"madrigal",
"london22",
"krakatoa",
"junction",
"intranet",
"humility",
"harmless",
"grace123",
"giuliana",
"gauntlet",
"fugitive",
"flatland",
"feelings",
"fabregas",
"emanuele",
"election",
"dumpster",
"douglas1",
"cruzeiro",
"cracking",
"control1",
"cheaters",
"centrino",
"captain1",
"canberra",
"botswana",
"atreides",
"asuncion",
"astroboy",
"aqualung",
"amnesiac",
"adorable",
"3edc4rfv",
"1z2x3c4v",
"19921992",
"14141414",
"12211221",
"yankees2",
"worldcup",
"vittorio",
"theworld",
"thebeast",
"thaddeus",
"telemark",
"sylvania",
"surveyor",
"suitcase",
"stroller",
"stripped",
"stallone",
"smoke420",
"septembe",
"sandberg",
"rousseau",
"revenant",
"pepsi123",
"pembroke",
"parkside",
"outbreak",
"obsolete",
"nutshell",
"nounours",
"nonenone",
"momentum",
"michele1",
"maldives",
"magdalen",
"lockhart",
"krokodil",
"humboldt",
"homebase",
"headshot",
"headless",
"hazelnut",
"gremlins",
"frankie1",
"frank123",
"fireman1",
"external",
"entering",
"dulcinea",
"dropkick",
"draconis",
"dont4get",
"domestic",
"darkwing",
"corporal",
"cocorico",
"chimaera",
"cheyanne",
"breakers",
"bluesman",
"bethesda",
"basketba",
"andyandy",
"allison1",
"Garfield",
"Abcd1234",
"yoyoyoyo",
"yeahbaby",
"wetpussy",
"variable",
"unicorn1",
"trillium",
"torrance",
"tikitiki",
"thumper1",
"thesaint",
"theforce",
"teiubesc",
"sweet123",
"succubus",
"stockman",
"steve123",
"speeding",
"sokrates",
"showboat",
"sequence",
"qwerty99",
"postcard",
"polkadot",
"orlando1",
"nicolas1",
"nicknick",
"naughty1",
"marielle",
"maneater",
"lionlion",
"leapfrog",
"kirkwood",
"kilkenny",
"jordan12",
"intercom",
"informix",
"hounddog",
"homicide",
"herschel",
"hatteras",
"harakiri",
"halfmoon",
"fivestar",
"firewood",
"executor",
"elcamino",
"egyptian",
"eclipse1",
"duckling",
"drumming",
"drifting",
"daisydog",
"coolgirl",
"contrast",
"choclate",
"chilling",
"channels",
"catapult",
"careless",
"californ",
"brendan1",
"beverley",
"atalanta",
"ashley12",
"arizona1",
"antihero",
"andrew12",
"allright",
"ab123456",
"43214321",
"18436572",
"windows7",
"wellcome",
"waldemar",
"valerian",
"tristan1",
"tornado1",
"thunders",
"tennyson",
"tarragon",
"tapestry",
"tajmahal",
"sunny123",
"struggle",
"starling",
"sobriety",
"snowfall",
"skyline1",
"shirley1",
"shalimar",
"settings",
"schnecke",
"satriani",
"sasha123",
"sailfish",
"roserose",
"qwerty22",
"prashant",
"powerman",
"powerade",
"plastics",
"pinkpink",
"parallel",
"papercut",
"p4ssword",
"navyseal",
"monopoli",
"mnemonic",
"millenia",
"membrane",
"manitoba",
"lineage2",
"leopards",
"karoline",
"johnpaul",
"interior",
"homepage",
"greeting",
"golfgolf",
"glassman",
"friction",
"filomena",
"ethereal",
"emotions",
"dudedude",
"douglass",
"dominika",
"demetrio",
"demented",
"decision",
"cuthbert",
"compound",
"comatose",
"civilwar",
"castello",
"cachorro",
"bulletin",
"brandnew",
"bluegill",
"baywatch",
"bastardo",
"bagheera",
"annalisa",
"allstate",
"alberto1",
"Samantha",
"78945612",
"01010101",
"yellow12",
"wildbill",
"whittier",
"vittoria",
"virgilio",
"trusting",
"troubles",
"tonytony",
"thebest1",
"terriers",
"template",
"telefoon",
"talented",
"supermen",
"starting",
"sixpence",
"sidewalk",
"shoshana",
"rainbow7",
"rafferty",
"qwerty77",
"qwerty00",
"pheasant",
"pentium3",
"patrizia",
"overlook",
"overhead",
"okokokok",
"nwo4life",
"novembre",
"newlife1",
"newdelhi",
"myspace1",
"myfriend",
"munchies",
"moneybag",
"molecule",
"mercury1",
"melville",
"mcintyre",
"mattress",
"maritime",
"mariachi",
"loveyou2",
"lovesong",
"lolalola",
"lindsey1",
"lifeboat",
"katie123",
"kasandra",
"jupiter1",
"julia123",
"india123",
"henry123",
"henrique",
"hardball",
"handbook",
"hacienda",
"grenoble",
"giuliano",
"freehand",
"fragment",
"foreskin",
"ensemble",
"eclectic",
"dogfight",
"dodgers1",
"diogenes",
"dillweed",
"demon666",
"daybreak",
"dagobert",
"culinary",
"crossing",
"controls",
"cobblers",
"charissa",
"buster12",
"bungalow",
"brianna1",
"bella123",
"ballroom",
"andre123",
"analysis",
"amber123",
"aa123456",
"2wsx3edc",
"12131213",
"wertwert",
"vivienne",
"tuppence",
"trafford",
"teddy123",
"streamer",
"star1234",
"sparrows",
"solomon1",
"sideshow",
"sherbert",
"sebastia",
"scribble",
"sarasota",
"sarasara",
"sarah123",
"sanguine",
"sandy123",
"robert12",
"redhorse",
"rational",
"radioman",
"qwerty01",
"poophead",
"phantoms",
"paperino",
"organize",
"optiplex",
"october1",
"neverdie",
"monsieur",
"monkfish",
"master01",
"marymary",
"lucas123",
"logistic",
"lemmings",
"langston",
"killer11",
"jack1234",
"ireland1",
"house123",
"hihihihi",
"hellhole",
"hardwood",
"funhouse",
"fiorella",
"farewell",
"fantasma",
"failsafe",
"explicit",
"esposito",
"duckduck",
"drilling",
"dragon10",
"dickweed",
"crunchie",
"crawfish",
"chessman",
"chanelle",
"chamonix",
"candy123",
"brainiac",
"birdland",
"binladen",
"billings",
"bareback",
"bacteria",
"asdfqwer",
"asd12345",
"arpeggio",
"anthony2",
"animator",
"amazonas",
"alpacino",
"adelaida",
"adamadam",
"aaron123",
"Einstein",
"90909090",
"1234zxcv",
"yamamoto",
"wormhole",
"whiteman",
"westgate",
"watchmen",
"vergeten",
"veracruz",
"vanquish",
"uuuuuuuu",
"trucking",
"trooper1",
"timelord",
"strangle",
"stoneman",
"starless",
"spagetti",
"sorensen",
"somethin",
"snowhite",
"slovakia",
"skydiver",
"silicone",
"silencio",
"selector",
"scramble",
"scott123",
"salinger",
"reminder",
"redheads",
"phaedrus",
"paulchen",
"passion1",
"paraguay",
"panda123",
"palacios",
"osbourne",
"onepiece",
"mutation",
"murakami",
"mercator",
"mario123",
"lynnette",
"lookatme",
"linda123",
"lightnin",
"lifeless",
"leopoldo",
"kristin1",
"knitting",
"katrina1",
"hershey1",
"gridlock",
"gigantic",
"fred1234",
"flatline",
"firehawk",
"fellatio",
"eruption",
"dragons1",
"dragon88",
"delorean",
"decipher",
"darkblue",
"creatine",
"counting",
"coolidge",
"cookie12",
"converge",
"clubbing",
"cbr600rr",
"carnegie",
"calabria",
"buttfuck",
"broncos1",
"blueball",
"beautifu",
"barnacle",
"babygurl",
"asturias",
"armchair",
"archives",
"aperture",
"amandine",
"22446688",
"20032003",
"19641964",
"12141214",
"01230123",
"yourname",
"warszawa",
"therock1",
"testuser",
"temp1234",
"swordfis",
"superdog",
"sunflowe",
"soccer22",
"slovenia",
"sinfonia",
"scimitar",
"rosebush",
"redriver",
"redeemed",
"ramstein",
"qweasdzx",
"plumbing",
"pickwick",
"parsifal",
"overcome",
"ninjutsu",
"newport1",
"newcomer",
"monkey01",
"minority",
"mariette",
"loveland",
"lagrange",
"kaitlynn",
"john1234",
"invictus",
"inventor",
"inspired",
"hurrican",
"honey123",
"holbrook",
"heracles",
"hathaway",
"governor",
"goodrich",
"gizmo123",
"friday13",
"fortytwo",
"foreplay",
"fishhook",
"fishfish",
"fillmore",
"espinoza",
"emerald1",
"edgewood",
"duisburg",
"drummers",
"dowjones",
"cameroon",
"buddyboy",
"bracelet",
"bogeyman",
"bluerose",
"birdcage",
"billy123",
"beepbeep",
"asdfgh12",
"antonina",
"anabolic",
"allister",
"albacore",
"airedale",
"activity",
"Patricia",
"99887766",
"20202020",
"19701970",
"yardbird",
"xcountry",
"wildrose",
"watanabe",
"wareagle",
"validate",
"tripping",
"treetree",
"timbuktu",
"summer00",
"stuntman",
"steelman",
"spartan1",
"snowshoe",
"smuggler",
"slowhand",
"shadow01",
"schuster",
"satelite",
"rightnow",
"r4e3w2q1",
"quagmire",
"porridge",
"peerless",
"paganini",
"optional",
"nowayout",
"newstart",
"neworder",
"monkey13",
"mission1",
"mcmillan",
"lucky777",
"lombardo",
"lindberg",
"larkspur",
"lambchop",
"lalaland",
"kirakira",
"joshua12",
"january1",
"infinito",
"identify",
"hellgate",
"heatwave",
"grounded",
"greenish",
"gorillaz",
"gerhardt",
"generous",
"gauthier",
"frontera",
"freezing",
"fracture",
"fastlane",
"drafting",
"donnelly",
"dolomite",
"damocles",
"critters",
"crickets",
"crabtree",
"cortland",
"comrades",
"clothing",
"checking",
"charmed1",
"cathleen",
"carter15",
"carleton",
"blueline",
"bigblack",
"bastard1",
"backspin",
"babababa",
"audition",
"argentum",
"antonius",
"antiques",
"abigail1",
"14531453",
"woodlawn",
"windward",
"warranty",
"visitors",
"trespass",
"trashcan",
"topnotch",
"tigger12",
"summer05",
"summer01",
"sturgeon",
"strikers",
"skipjack",
"shipyard",
"shekinah",
"scouting",
"sanpedro",
"sandrock",
"rootroot",
"ronaldo9",
"reynaldo",
"relative",
"radagast",
"qwertzui",
"presidio",
"presence",
"prentice",
"playback",
"philippa",
"peterman",
"peregrin",
"peaceman",
"papabear",
"organist",
"octavian",
"nascar24",
"monteiro",
"monkeys1",
"metaphor",
"manifold",
"makelove",
"lysander",
"lobsters",
"julie123",
"johngalt",
"jamaica1",
"jalapeno",
"jacobsen",
"isengard",
"hutchins",
"horizons",
"hawkwind",
"happyboy",
"gutentag",
"gracious",
"glenwood",
"frogfrog",
"fraction",
"folklore",
"fantasy1",
"express1",
"exposure",
"everton1",
"employee",
"economic",
"ducksoup",
"diskette",
"delacruz",
"creepers",
"clements",
"cheerful",
"catering",
"capucine",
"capacity",
"bridgett",
"boyscout",
"bingo123",
"belgrade",
"beginner",
"bavarian",
"backfire",
"astaroth",
"arsehole",
"annelise",
"andrew01",
"anabelle",
"albright",
"airlines",
"adelante",
"account1",
"Maverick",
"85208520",
"14121412",
"yahoo123",
"wretched",
"winthrop",
"westwind",
"weinberg",
"trashman",
"toronto1",
"thomas01",
"thibault",
"syndrome",
"swinging",
"sweetest",
"sunburst",
"sperling",
"spectral",
"soldier1",
"silmaril",
"shoulder",
"shahrukh",
"settlers",
"scotsman",
"scofield",
"schumann",
"rockrock",
"rockland",
"qwerty69",
"promises",
"priscila",
"priority",
"playoffs",
"pebbles1",
"overseer",
"opposite",
"octavius",
"nikenike",
"nehemiah",
"mystery1",
"morticia",
"monkey11",
"misty123",
"milenium",
"michael3",
"lincoln1",
"lilwayne",
"lausanne",
"kokokoko",
"kilowatt",
"jacob123",
"interval",
"ignorant",
"huntsman",
"homesick",
"highbury",
"hellbent",
"guerilla",
"graywolf",
"grandson",
"gargamel",
"gameplay",
"firefly1",
"fighter1",
"fielding",
"familiar",
"falconer",
"ezequiel",
"dynamics",
"demetria",
"darkroom",
"curtains",
"currency",
"crocodil",
"crawling",
"christy1",
"chivalry",
"charlie7",
"catriona",
"carolann",
"cantona7",
"canfield",
"buttocks",
"brinkley",
"bordello",
"blissful",
"blackbox",
"billiard",
"bigbooty",
"bastille",
"as123456",
"artofwar",
"annalena",
"animated",
"alvarado",
"alicante",
"alex2000",
"accurate",
"17171717",
"123456as",
"00112233",
"password",
"12345678",
"1q2w3e4r",
"sunshine",
"football",
"computer",
"superman",
"internet",
"iloveyou",
"1qaz2wsx",
"baseball",
"whatever",
"princess",
"abcd1234",
"starwars",
"trustno1",
"jennifer",
"michelle",
"mercedes",
"benjamin",
"11111111",
"samantha",
"victoria",
"asdf1234",
"1234qwer",
"q1w2e3r4",
"elephant",
"garfield",
"jonathan",
"caroline",
"maverick",
"midnight",
"88888888",
"creative",
"cocacola",
"passw0rd",
"blink182",
"danielle",
"scorpion",
"veronica",
"nicholas",
"asdfasdf",
"december",
"patricia",
"security",
"slipknot",
"november",
"jordan23",
"qwertyui",
"carolina",
"hardcore",
"corvette",
"12341234",
"remember",
"qwer1234",
"leonardo",
"snickers",
"williams",
"angelina",
"anderson",
"pakistan",
"marlboro",
"kimberly",
"00000000",
"snowball",
"godzilla",
"hello123",
"champion",
"precious",
"einstein",
"napoleon",
"mountain",
"dolphins",
"fernando",
"87654321",
"paradise",
"motorola",
"bullshit",
"brooklyn",
"qwerty12",
"franklin",
"american",
"platinum",
"icecream",
"darkness",
"cristina",
"colorado",
"steelers",
"serenity",
"mitchell",
"lollipop",
"marshall",
"1qazxsw2",
"12344321",
"startrek",
"business",
"nintendo",
"12qwaszx",
"asdfghjk",
"Password",
"zaq12wsx",
"scotland",
"hercules",
"explorer",
"firebird",
"engineer",
"virginia",
"simpsons",
"angelica",
"isabelle",
"isabella",
"changeme",
"passport",
"infinity",
"courtney",
"scarface",
"pavilion",
"abcdefgh",
"a1b2c3d4",
"harrison",
"spitfire",
"birthday",
"guinness",
"logitech",
"emmanuel",
"11223344",
"goldfish",
"cheyenne",
"testtest",
"stargate",
"anything",
"aaaaaaaa",
"welcome1",
"eternity",
"westside",
"maryjane",
"michael1",
"lawrence",
"kristina",
"kawasaki",
"drowssap",
"blahblah",
"babygirl",
"poohbear",
"florence",
"sapphire",
"hamilton",
"greenday",
"twilight",
"swimming",
"stardust",
"predator",
"penelope",
"michigan",
"margaret",
"brittany",
"shithead",
"redskins",
"pussycat",
"fireball",
"cherokee",
"1234abcd",
"lovelove",
"thailand",
"lasvegas",
"butthead",
"blizzard",
"shamrock",
"bluebird",
"atlantis",
"magnolia",
"juventus",
"diamonds",
"warcraft",
"renegade",
"mohammed",
"shopping",
"savannah",
"giovanni",
"12121212",
"wildcats",
"portugal",
"santiago",
"kathleen",
"clifford",
"55555555",
"rosemary",
"vacation",
"chandler",
"99999999",
"lorraine",
"children",
"beatrice",
"airborne",
"valentin",
"kamikaze",
"software",
"22222222",
"salvador",
"panthers",
"lacrosse",
"charlie1",
"cardinal",
"bluemoon",
"zeppelin",
"rockstar",
"operator",
"dickhead",
"anaconda",
"77777777",
"skittles",
"personal",
"kingkong",
"geronimo",
"robinson",
"kingston",
"hannibal",
"download",
"darkstar",
"sweetpea",
"softball",
"pa55word",
"keyboard",
"darkside",
"assassin",
"vladimir",
"national",
"matthew1",
"brothers",
"warriors",
"universe",
"rush2112",
"mushroom",
"bigdaddy",
"1a2b3c4d",
"ultimate",
"peterpan",
"loverboy",
"truelove",
"trombone",
"madeline",
"gangster",
"dingdong",
"catalina",
"kittycat",
"aquarius",
"patriots",
"ihateyou",
"blessing",
"airplane",
"stingray",
"hellfire",
"guardian",
"flamingo",
"socrates",
"richmond",
"electric",
"thankyou",
"sterling",
"munchkin",
"morpheus",
"imperial",
"goodluck",
"columbia",
"campbell",
"oblivion",
"freedom1",
"valencia",
"spectrum",
"jessica1",
"jeremiah",
"handsome",
"goldberg",
"gabriela",
"anthony1",
"a1234567",
"xxxxxxxx",
"peekaboo",
"montreal",
"kangaroo",
"immortal",
"chocolat",
"thompson",
"research",
"oklahoma",
"mariposa",
"defender",
"applepie",
"squirrel",
"hongkong",
"dinosaur",
"babydoll",
"wolfgang",
"semperfi",
"patience",
"fletcher",
"drpepper",
"creation",
"wordpass",
"passwort",
"original",
"martinez",
"labrador",
"apple123",
"sundance",
"redwings",
"monopoly",
"lionking",
"director",
"44444444",
"sherlock",
"marianne",
"lancelot",
"jeanette",
"cannabis",
"werewolf",
"marathon",
"longhorn",
"happy123",
"brucelee",
"wrangler",
"william1",
"stranger",
"scarlett",
"morrison",
"february",
"fantasia",
"designer",
"bulldogs",
"sullivan",
"saturday",
"pingpong",
"kristine",
"fuckyou1",
"fearless",
"airforce",
"theodore",
"starfish",
"pass1234",
"cinnamon",
"overlord",
"michaela",
"meredith",
"abc12345",
"aardvark",
"Passw0rd",
"trinidad",
"thursday",
"standard",
"pearljam",
"springer",
"ragnarok",
"portland",
"nathalie",
"lemonade",
"lavender",
"gotohell",
"freckles",
"crusader",
"commando",
"clarence",
"cadillac",
"verbatim",
"umbrella",
"splinter",
"register",
"qwert123",
"penguins",
"ncc1701d",
"estrella",
"downtown",
"colombia",
"bollocks",
"69696969",
"showtime",
"qwerasdf",
"mongoose",
"illusion",
"cooldude",
"treasure",
"monalisa",
"justdoit",
"ericsson",
"chelsea1",
"achilles",
"a1s2d3f4",
"veronika",
"test1234",
"sporting",
"papillon",
"juliette",
"fuckyou2",
"firewall",
"cristian",
"cavalier",
"canadian",
"admin123",
"together",
"pa55w0rd",
"halflife",
"formula1",
"thirteen",
"rastaman",
"mustang1",
"cucumber",
"sheridan",
"qqqqqqqq",
"punisher",
"lovelife",
"gretchen",
"chevelle",
"chester1",
"wireless",
"sandiego",
"pokemon1",
"lollypop",
"gorgeous",
"chickens",
"blackman",
"atlantic",
"wildfire",
"waterloo",
"james123",
"homework",
"highland",
"eldorado",
"discover",
"alphabet",
"zaq1xsw2",
"tropical",
"question",
"presario",
"notebook",
"nebraska",
"bullseye",
"valhalla",
"tomorrow",
"richard1",
"positive",
"plymouth",
"patrick1",
"faithful",
"doberman",
"criminal",
"crackers",
"converse",
"casanova",
"attitude",
"66666666",
"scooter1",
"rochelle",
"punkrock",
"kentucky",
"insomnia",
"hooligan",
"gertrude",
"blueeyes",
"terminal",
"poseidon",
"paranoid",
"laurence",
"istanbul",
"frederic",
"doomsday",
"bradford",
"bonehead",
"apollo13",
"westwood",
"satan666",
"reynolds",
"mckenzie",
"magician",
"innocent",
"hotstuff",
"fountain",
"concrete",
"capslock",
"snuggles",
"megadeth",
"medicine",
"jackson1",
"intrepid",
"green123",
"geoffrey",
"dynamite",
"columbus",
"chemical",
"chargers",
"username",
"sherwood",
"moonbeam",
"meowmeow",
"matthias",
"jackson5",
"honolulu",
"diamond1",
"crawford",
"broadway",
"zzzzzzzz",
"whocares",
"svetlana",
"southern",
"pleasure",
"makaveli",
"honeybee",
"francois",
"chicken1",
"bookworm",
"PASSWORD",
"33333333",
"sunlight",
"stallion",
"katerina",
"hedgehog",
"happyday",
"davidson",
"cerberus",
"blackcat",
"arsenal1",
"angel123",
"10101010",
"training",
"republic",
"recovery",
"maradona",
"intruder",
"hermione",
"hastings",
"goldstar",
"fredfred",
"federico",
"deftones",
"blackout",
"1234567a",
"wolfpack",
"thunder1",
"tacobell",
"solution",
"shanghai",
"rootbeer",
"phillips",
"monsters",
"lonewolf",
"keystone",
"johannes",
"grateful",
"continue",
"confused",
"brighton",
"yankees1",
"triangle",
"peterson",
"marianna",
"mandrake",
"inuyasha",
"hardware",
"freebird",
"ferguson",
"dominick",
"bullfrog",
"babylon5",
"13131313",
"zanzibar",
"transfer",
"sparkles",
"shepherd",
"resident",
"property",
"pictures",
"mischief",
"kristian",
"heineken",
"hahahaha",
"eastside",
"daffodil",
"charming",
"billybob",
"adelaide",
"underdog",
"technics",
"samsung1",
"phoenix1",
"musicman",
"marjorie",
"letmein1",
"hospital",
"handball",
"gonzales",
"budapest",
"brandon1",
"alliance",
"adrienne",
"aberdeen",
"thuglife",
"sentinel",
"richards",
"newyork1",
"mortimer",
"marcello",
"magazine",
"infantry",
"hopeless",
"fandango",
"deadhead",
"clarissa",
"christie",
"charlene",
"billyboy",
"bangbang",
"absolute",
"titanium",
"tiger123",
"superior",
"stefanie",
"spaceman",
"somebody",
"sinclair",
"pppppppp",
"mmmmmmmm",
"military",
"loveless",
"karolina",
"fernanda",
"felicity",
"dietcoke",
"brewster",
"babyblue",
"ashleigh",
"14789632",
"whiskers",
"valkyrie",
"superfly",
"strength",
"progress",
"muhammad",
"maryland",
"daughter",
"clarinet",
"chuckles",
"almighty",
"1qaz1qaz",
"sneakers",
"saratoga",
"qawsedrf",
"majestic",
"kingfish",
"japanese",
"graphics",
"flounder",
"coltrane",
"chris123",
"checkers",
"barbados",
"augustus",
"angelika",
"washburn",
"survivor",
"stanford",
"soulmate",
"rasputin",
"pallmall",
"overkill",
"meatloaf",
"lowrider",
"katarina",
"ilovegod",
"heather1",
"hallo123",
"giuseppe",
"eastwood",
"dominion",
"chiquita",
"chipmunk",
"castillo",
"berkeley",
"thinking",
"tarheels",
"seminole",
"pornstar",
"platypus",
"nirvana1",
"mephisto",
"johnjohn",
"gameover",
"fuckface",
"david123",
"darklord",
"cutiepie",
"carnival",
"candyman",
"blowfish",
"ssssssss",
"sandwich",
"sailboat",
"mandarin",
"knuckles",
"jasmine1",
"hardrock",
"boomboom",
"benedict",
"babyface",
"albatros",
"sprinter",
"rolltide",
"r2d2c3po",
"mustangs",
"missouri",
"meridian",
"meatball",
"malaysia",
"killbill",
"illinois",
"gonzalez",
"georgina",
"gargoyle",
"disaster",
"complete",
"claymore",
"chainsaw",
"bluebell",
"98765432",
"wishbone",
"vampires",
"smashing",
"rhiannon",
"rachelle",
"playtime",
"marcella",
"lonestar",
"heritage",
"hayabusa",
"forsaken",
"ferrari1",
"backdoor",
"asshole1",
"11235813",
"yosemite",
"yogibear",
"talisman",
"syracuse",
"randolph",
"raistlin",
"preacher",
"millions",
"metallic",
"madison1",
"dontknow",
"coolcool",
"charisma",
"sinister",
"passpass",
"mohammad",
"mcdonald",
"frontier",
"flipflop",
"eggplant",
"dannyboy",
"daniella",
"chrysler",
"cameron1",
"buckshot",
"arkansas",
"america1",
"12345679",
"romantic",
"robotics",
"redalert",
"megatron",
"mamapapa",
"hyperion",
"gabriel1",
"fuckfuck",
"friendly",
"florida1",
"dreaming",
"doghouse",
"christin",
"brigitte",
"addicted",
"shadow12",
"porkchop",
"negative",
"mistress",
"melissa1",
"jermaine",
"james007",
"francine",
"delphine",
"crystal1",
"chestnut",
"auckland",
"wanderer",
"tomahawk",
"thanatos",
"snoopdog",
"roderick",
"princesa",
"pentagon",
"money123",
"mechanic",
"creature",
"cornwall",
"chadwick",
"calendar",
"abdullah",
"vendetta",
"stephane",
"revolver",
"railroad",
"p4ssw0rd",
"mariners",
"holyshit",
"database",
"bobafett",
"bernardo",
"amethyst",
"advanced",
"whistler",
"slamdunk",
"scrabble",
"roadkill",
"rainbows",
"polopolo",
"obsidian",
"northern",
"learning",
"elements",
"electron",
"customer",
"brisbane",
"baritone",
"amarillo",
"alexandr",
"12301230",
"windmill",
"vanhalen",
"surprise",
"starfire",
"speakers",
"ncc1701e",
"lifetime",
"kittykat",
"fredrick",
"fidelity",
"fabulous",
"everyday",
"coolness",
"concorde",
"catwoman",
"babybaby",
"vodafone",
"traveler",
"rainbow1",
"potatoes",
"pipeline",
"philippe",
"monterey",
"lipstick",
"lakeside",
"insanity",
"fishbone",
"bordeaux",
"21122112",
"windsurf",
"velocity",
"vagabond",
"reloaded",
"raindrop",
"prudence",
"pharmacy",
"peaceful",
"marietta",
"letmein2",
"ladybird",
"internal",
"gigabyte",
"fourteen",
"dolphin1",
"chambers",
"bunghole",
"buckeyes",
"bluefish",
"23232323",
"12369874",
"zerocool",
"wrestler",
"tortoise",
"sysadmin",
"starship",
"qwerty11",
"primrose",
"politics",
"paranoia",
"pancakes",
"overload",
"matthews",
"marriage",
"macaroni",
"jonathon",
"jackjack",
"infinite",
"heinrich",
"graduate",
"goodness",
"godspeed",
"feedback",
"cornelia",
"corleone",
"choochoo",
"chairman",
"butthole",
"buddy123",
"azsxdcfv",
"sleeping",
"pringles",
"power123",
"paradigm",
"nickolas",
"nautilus",
"feathers",
"facebook",
"dragon12",
"brittney",
"aviation",
"19841984",
"10203040",
"wildwood",
"thrasher",
"speedway",
"songbird",
"sickness",
"shannon1",
"screamer",
"monster1",
"mauricio",
"love1234",
"devil666",
"budlight",
"ambrosia",
"adrianna",
"zxcvbnm1",
"windows1",
"toulouse",
"tazmania",
"slapshot",
"ministry",
"mathilde",
"lighting",
"helsinki",
"gateway1",
"fussball",
"frederik",
"flexible",
"festival",
"destiny1",
"daydream",
"coventry",
"constant",
"charles1",
"angeline",
"woodland",
"skinhead",
"sandrine",
"rockford",
"merchant",
"greatest",
"everlast",
"espresso",
"elizabet",
"dddddddd",
"chouchou",
"charlton",
"carlitos",
"blueblue",
"awesome1",
"aspirine",
"12345abc",
"stronger",
"starbuck",
"skeleton",
"scissors",
"reginald",
"redeemer",
"normandy",
"luckydog",
"laserjet",
"just4fun",
"greenbay",
"graffiti",
"doughboy",
"dortmund",
"building",
"bbbbbbbb",
"annabell",
"zimbabwe",
"tunafish",
"thisisit",
"stafford",
"spalding",
"solitude",
"robotech",
"rainbow6",
"qazwsx12",
"pooppoop",
"minister",
"leonidas",
"kirkland",
"integral",
"ilovesex",
"ignatius",
"heavenly",
"gggggggg",
"exchange",
"bulldog1",
"blackdog",
"bearbear",
"winfield",
"westlife",
"thriller",
"spartans",
"sausages",
"printing",
"palmtree",
"opendoor",
"mosquito",
"milkyway",
"laughter",
"klondike",
"kingsley",
"jesus123",
"humphrey",
"hillside",
"hattrick",
"function",
"fighting",
"delaware",
"costello",
"catalyst",
"babylove",
"assholes",
"andersen",
"alexande",
"19891989",
"1234asdf",
"whiplash",
"tiffany1",
"sammy123",
"rockwell",
"reddevil",
"maxwell1",
"gordon24",
"glendale",
"giovanna",
"foxylady",
"fortress",
"favorite",
"doughnut",
"comanche",
"cheshire",
"cherries",
"catarina",
"bertrand",
"barefoot",
"arabella",
"vanguard",
"stephen1",
"rhapsody",
"reckless",
"pumpkin1",
"powerful",
"painting",
"nocturne",
"nickname",
"mynameis",
"mikemike",
"llllllll",
"leighton",
"kkkkkkkk",
"johnston",
"holidays",
"handyman",
"fuckoff1",
"front242",
"flamenco",
"escalade",
"division",
"covenant",
"cannibal",
"annmarie",
"alcatraz",
"11112222",
"wwwwwwww",
"wildcard",
"whitesox",
"vincent1",
"thornton",
"survival",
"sprocket",
"somerset",
"skorpion",
"services",
"restless",
"pumpkins",
"meathead",
"lucky123",
"licorice",
"language",
"jackass1",
"infiniti",
"gamecube",
"flanders",
"disciple",
"diplomat",
"crescent",
"catholic",
"capoeira",
"browning",
"biscuits",
"alexalex",
"P@ssw0rd",
"Jennifer",
"19861986",
"winston1",
"violator",
"super123",
"straight",
"sorcerer",
"sidekick",
"shredder",
"schubert",
"prestige",
"peter123",
"nonsense",
"mulligan",
"moneyman",
"matchbox",
"marauder",
"longhair",
"lisalisa",
"kayleigh",
"islander",
"genesis1",
"gardenia",
"gabriele",
"edmonton",
"downhill",
"digital1",
"cromwell",
"chowchow",
"carebear",
"vanessa1",
"terrapin",
"stockton",
"smoothie",
"seahawks",
"rebecca1",
"rangers1",
"puppydog",
"marigold",
"gregorio",
"gangbang",
"dutchess",
"daylight",
"clueless",
"calamity",
"beefcake",
"aquarium",
"anathema",
"ambition",
"19821982",
"wildlife",
"snowbird",
"qwerqwer",
"prospect",
"natalie1",
"lockdown",
"italiano",
"irishman",
"infamous",
"hydrogen",
"hartford",
"goodyear",
"generals",
"garrison",
"foxhound",
"entrance",
"eighteen",
"diamante",
"daedalus",
"cocktail",
"caligula",
"borabora",
"behemoth",
"balloons",
"bachelor",
"waterman",
"teenager",
"spanking",
"soccer10",
"sergeant",
"seashell",
"seahorse",
"riffraff",
"possible",
"pinnacle",
"nostromo",
"latitude",
"kevin123",
"invasion",
"hibiscus",
"hallmark",
"envision",
"charcoal",
"blue1234",
"antelope",
"aircraft",
"123456aa",
"viktoria",
"stripper",
"stefania",
"smirnoff",
"seraphim",
"ronaldo7",
"reporter",
"raiders1",
"nineteen",
"monolith",
"memories",
"memorial",
"massacre",
"honduras",
"goofball",
"fullmoon",
"forever1",
"elefante",
"doorknob",
"dipstick",
"commerce",
"carousel",
"callisto",
"berenice",
"asdfzxcv",
"alex1234",
"Welcome1",
"19871987",
"wormwood",
"starstar",
"sexygirl",
"rosewood",
"roadster",
"rapunzel",
"prisoner",
"prescott",
"pizza123",
"phillies",
"phantom1",
"perfect1",
"pasadena",
"optimist",
"master12",
"junkmail",
"inspiron",
"hhhhhhhh",
"griffith",
"golfball",
"forester",
"euphoria",
"england1",
"death666",
"conquest",
"clitoris",
"cartoons",
"buckaroo",
"bluejays",
"violence",
"testpass",
"terrence",
"temporal",
"teamwork",
"spencer1",
"shipping",
"roosters",
"prophecy",
"popcorn1",
"playmate",
"panorama",
"p0o9i8u7",
"landmark",
"johnson1",
"iverson3",
"instinct",
"infected",
"honeydew",
"document",
"deadline",
"cowboys1",
"climbing",
"bubbles1",
"bluestar",
"bathroom",
"anamaria",
"25802580",
"24682468",
"whiteboy",
"titleist",
"tiberius",
"retarded",
"palomino",
"outsider",
"oooooooo",
"musician",
"michelin",
"hyacinth",
"gatorade",
"fuzzball",
"everyone",
"delirium",
"daisy123",
"critical",
"cordelia",
"capitals",
"caliente",
"bobdylan",
"Michelle",
"1a2s3d4f",
"19781978",
"voltaire",
"thedoors",
"special1",
"southpaw",
"soccer12",
"ruthless",
"reaction",
"qazwsxed",
"portable",
"passcode",
"official",
"mindless",
"masamune",
"lalalala",
"holloway",
"hairball",
"dirtbike",
"dilligaf",
"clippers",
"chicago1",
"caldwell",
"agent007",
"19831983",
"19801980",
"19751975",
"warrior1",
"vertical",
"timeless",
"thegreat",
"spelling",
"slippery",
"rrrrrrrr",
"ricochet",
"protocol",
"producer",
"penguin1",
"p455w0rd",
"olivetti",
"oliveira",
"metalica",
"mannheim",
"mandingo",
"magellan",
"machines",
"lovebird",
"jason123",
"inflames",
"headache",
"godbless",
"gemstone",
"ffffffff",
"cyclones",
"colonial",
"claudius",
"bulgaria",
"brunette",
"bradshaw",
"bastards",
"basement",
"acapulco",
"25252525",
"12312312",
"zachary1",
"yingyang",
"workshop",
"trueblue",
"sycamore",
"stigmata",
"sabrina1",
"riccardo",
"playboy1",
"override",
"music123",
"mortgage",
"meandyou",
"macdaddy",
"knockers",
"kisskiss",
"jjjjjjjj",
"hysteria",
"forgiven",
"distance",
"cosworth",
"coconuts",
"carlisle",
"asdfjkl;",
"31415926",
"21212121",
"yokohama",
"tommy123",
"sheepdog",
"seinfeld",
"sabotage",
"pressure",
"pinetree",
"pavement",
"oriental",
"offshore",
"netscape",
"michaels",
"mash4077",
"mallorca",
"junkyard",
"johncena",
"jakejake",
"hawthorn",
"hawaiian",
"frenchie",
"fishing1",
"fastball",
"deathrow",
"calimero",
"breakout",
"black123",
"bismarck",
"alkaline",
"zxcv1234",
"tryagain",
"thatcher",
"stampede",
"scheisse",
"sayonara",
"passions",
"nothing1",
"nameless",
"mysterio",
"monkey12",
"millwall",
"megabyte",
"mccarthy",
"magister",
"madhouse",
"liverpoo",
"laetitia",
"jennings",
"holstein",
"freefall",
"flawless",
"ebenezer",
"divinity",
"delpiero",
"chastity",
"charlott",
"carlotta",
"buchanan",
"bradley1",
"aventura",
"asdffdsa",
"19741974",
"zildjian",
"wargames",
"vvvvvvvv",
"unicorns",
"tenerife",
"tasmania",
"symphony",
"splendid",
"sonyvaio",
"snapshot",
"saunders",
"sarajevo",
"reverend",
"polaroid",
"perfecto",
"nokia123",
"natasha1",
"mystical",
"melanie1",
"material",
"maddison",
"landlord",
"juvenile",
"goodwill",
"goldwing",
"gilberto",
"gandalf1",
"fuckthis",
"flapjack",
"flamengo",
"finnegan",
"fabienne",
"erection",
"clemente",
"caterina",
"capetown",
"antonio1",
"angelito",
"accounts",
"abstract",
"19911991",
"19761976",
"01234567",
"vincenzo",
"townsend",
"soccer11",
"smithers",
"shooting",
"shitshit",
"senators",
"redbaron",
"percival",
"painless",
"myfamily",
"mongolia",
"miroslav",
"macarena",
"lakewood",
"killer12",
"incoming",
"immanuel",
"hometown",
"homeless",
"giordano",
"genocide",
"enforcer",
"dispatch",
"codename",
"cccccccc",
"caramelo",
"callaway",
"calculus",
"brian123",
"blessed1",
"attorney",
"asteroid",
"academia",
"12131415",
"yamahar1",
"tricolor",
"terrance",
"summer99",
"stirling",
"stamford",
"stairway",
"soldiers",
"shitface",
"scorpio1",
"principe",
"pizzahut",
"patricio",
"passwerd",
"mulberry",
"luscious",
"lifeline",
"legoland",
"kickflip",
"kennwort",
"kathrine",
"josefina",
"jesus777",
"hellsing",
"drummond",
"delldell",
"cupcakes",
"claudine",
"ciaociao",
"christia",
"cashmere",
"carthage",
"bookmark",
"bartlett",
"alphonse",
"Benjamin",
"51505150",
"woodside",
"vaseline",
"trinity1",
"toxicity",
"tommyboy",
"ticktock",
"teachers",
"strategy",
"stephens",
"snowdrop",
"smeghead",
"shutdown",
"sexysexy",
"popsicle",
"petersen",
"oscar123",
"maryanne",
"magicman",
"kingking",
"identity",
"icehouse",
"hannover",
"glorious",
"forgetit",
"fishtank",
"epiphone",
"elevator",
"elegance",
"drumline",
"devilman",
"delivery",
"chrissie",
"carnaval",
"caffeine",
"bukowski",
"brownies",
"bearcats",
"akatsuki",
"19941994",
"woofwoof",
"virginie",
"untitled",
"tttttttt",
"timothy1",
"stickman",
"starlite",
"smarties",
"oxymoron",
"oleander",
"ncc1701a",
"muhammed",
"morphine",
"mobydick",
"meltdown",
"medieval",
"mahogany",
"magic123",
"longshot",
"lockheed",
"livewire",
"lakeland",
"kenworth",
"interpol",
"hunter12",
"hibernia",
"helpdesk",
"godofwar",
"fishhead",
"ethernet",
"duracell",
"crystals",
"colossus",
"besiktas",
"backlash",
"academic",
"abnormal",
"19901990",
"violetta",
"vineyard",
"terrible",
"suburban",
"stocking",
"snuffles",
"sideways",
"schwartz",
"salasana",
"rosalind",
"purchase",
"practice",
"poiuytre",
"piramide",
"montrose",
"molly123",
"maximus1",
"mammamia",
"lunchbox",
"lonesome",
"limerick",
"liberty1",
"ignition",
"homebrew",
"harry123",
"greenman",
"godsmack",
"firefire",
"daniel12",
"cricket1",
"contract",
"conflict",
"comeback",
"coldplay",
"believer",
"beaumont",
"angelita",
"23456789",
"woodward",
"wolverin",
"wellness",
"swingers",
"solstice",
"scratchy",
"rockport",
"redlight",
"puppy123",
"paulette",
"panther1",
"overtime",
"nazareth",
"mudvayne",
"movement",
"miracles",
"mike1234",
"maserati",
"marbella",
"kiwikiwi",
"jurassic",
"infernal",
"hereford",
"goodtime",
"goodlife",
"goodgirl",
"gamecock",
"gabriell",
"friends1",
"ferreira",
"ethiopia",
"dionysus",
"deadpool",
"christos",
"chauncey",
"castaway",
"carefree",
"burnside",
"borussia",
"bohemian",
"blackice",
"bigmouth",
"baptiste",
"augustin",
"asdfg123",
"alistair",
"advocate",
"adgjmptw",
"acoustic",
"Princess",
"19811981",
"11221122",
"youandme",
"vinicius",
"vauxhall",
"tyler123",
"terminus",
"surround",
"soccer13",
"sexylady",
"sessions",
"scirocco",
"schiller",
"schedule",
"rosebud1",
"regional",
"radiance",
"pioneers",
"phantasy",
"peaches1",
"p@ssw0rd",
"neutrino",
"kendrick",
"hogwarts",
"heinlein",
"guitarra",
"gillette",
"germania",
"flowers1",
"fighters",
"fastback",
"fabrizio",
"exercise",
"envelope",
"element1",
"eeeeeeee",
"doraemon",
"diabetes",
"damascus",
"coronado",
"cashflow",
"cardigan",
"blackboy",
"bitchass",
"backpack",
"anakonda",
"Victoria",
"911turbo",
"19851985",
"19721972",
"water123",
"viscount",
"violette",
"undertow",
"teacher1",
"success1",
"stephani",
"redstone",
"premiere",
"planning",
"paramore",
"packers1",
"nitrogen",
"natascha",
"moonwalk",
"maurizio",
"marzipan",
"mandolin",
"mamamama",
"maintain",
"macgyver",
"ludacris",
"loredana",
"killkill",
"justice1",
"jailbird",
"goodnews",
"freshman",
"firestar",
"eleonora",
"dragon11",
"domenico",
"discreet",
"crossbow",
"choppers",
"betrayed",
"bernhard",
"basilisk",
"antigone",
"alterego",
"alhambra",
"aerobics",
"Superman",
"20012001",
"1million",
"yyyyyyyy",
"woodruff",
"vampire1",
"tequiero",
"sunnyboy",
"specialk",
"sorrento",
"reliance",
"q2w3e4r5",
"proverbs",
"playgirl",
"pentium4",
"pedigree",
"partners",
"orange12",
"observer",
"nnnnnnnn",
"newworld",
"moriarty",
"minotaur",
"location",
"knockout",
"knickers",
"jeffrey1",
"hellyeah",
"greentea",
"goodgood",
"germany1",
"gasoline",
"flashman",
"fatality",
"emiliano",
"ellipsis",
"disorder",
"deadlock",
"davidoff",
"couscous",
"congress",
"cleaning",
"clarkson",
"charlie2",
"ceramics",
"casandra",
"cambodia",
"bigmoney",
"backbone",
"74108520",
"24681012",
"24242424",
"19881988",
"whatwhat",
"watching",
"tomatoes",
"tiramisu",
"tiberian",
"thurston",
"spinning",
"slippers",
"simon123",
"response",
"reindeer",
"porsche1",
"panchito",
"montana1",
"mayfield",
"marquise",
"manifest",
"magnetic",
"lovelace",
"lesbians",
"joystick",
"industry",
"gulliver",
"ganymede",
"galactic",
"esoteric",
"dropdead",
"drinking",
"devildog",
"copeland",
"christop",
"cheerios",
"chatting",
"changeit",
"cerulean",
"cabernet",
"bionicle",
"baltazar",
"amoremio",
"alpha123",
"alleycat",
"accident",
"19771977",
"123mudar",
"tingting",
"thething",
"testing1",
"tallulah",
"symmetry",
"summer69",
"smartass",
"shadow11",
"salesman",
"rushmore",
"resource",
"pregnant",
"pleasant",
"plankton",
"pendulum",
"paterson",
"partizan",
"olympics",
"networks",
"mystique",
"mckinley",
"mcgregor",
"maxpower",
"livelife",
"kokakola",
"katherin",
"julianna",
"jeannine",
"horseman",
"homeland",
"holiday1",
"hennessy",
"guesswho",
"greywolf",
"gilligan",
"gallardo",
"freewill",
"francis1",
"fordf150",
"fantomas",
"dutchman",
"drummer1",
"dementia",
"berliner",
"20002000",
"19951995",
"woodwork",
"winifred",
"welcome2",
"waterboy",
"troopers",
"theodora",
"sometime",
"russell1",
"roadking",
"rifleman",
"raymond1",
"qwerty13",
"priyanka",
"private1",
"pizzaman",
"phantasm",
"pathetic",
"nicotine",
"mollydog",
"minstrel",
"matthieu",
"maria123",
"lebron23",
"lakers24",
"kitty123",
"kindness",
"hatfield",
"getmoney",
"general1",
"forsythe",
"fontaine",
"feelgood",
"evidence",
"erickson",
"enter123",
"downfall",
"deadwood",
"crazyman",
"citation",
"calliope",
"broccoli",
"bleeding",
"bergkamp",
"asmodeus",
"artistic",
"antilles",
"anteater",
"anhyeuem",
"aaaa1111",
"Sunshine",
"Jonathan",
"19731973",
"19691969",
"wrinkles",
"trumpet1",
"triplets",
"sunnyday",
"summer12",
"students",
"start123",
"sopranos",
"siberian",
"shetland",
"sheppard",
"scrapper",
"schooner",
"pershing",
"parasite",
"pantera1",
"palmetto",
"overture",
"odysseus",
"noisette",
"narayana",
"nakamura",
"mediator",
"mcintosh",
"mazda626",
"marykate",
"manpower",
"malamute",
"justin12",
"jeronimo",
"jeremias",
"jamaican",
"imperium",
"humberto",
"hotmail1",
"hoosiers",
"goldmine",
"futurama",
"elisabet",
"dumpling",
"dragster",
"dragon13",
"dominica",
"dominate",
"dictator",
"cookbook",
"concerto",
"christel",
"beholder",
"babushka",
"autobahn",
"anywhere",
"acidburn",
"abhishek",
"z1x2c3v4",
"whiteout",
"topolino",
"thousand",
"thorsten",
"symantec",
"stanley1",
"splatter",
"sonysony",
"schaefer",
"reddwarf",
"position",
"popopopo",
"pikapika",
"piercing",
"pasquale",
"neighbor",
"mireille",
"lovesick",
"loverman",
"london12",
"lockwood",
"kowalski",
"kerberos",
"kellyann",
"jimmy123",
"jayhawks",
"innuendo",
"ilovemom",
"iiiiiiii",
"houston1",
"horrible",
"himalaya",
"highlife",
"hetfield",
"graphite",
"funnyman",
"f00tball",
"epiphany",
"elvis123",
"discount",
"danny123",
"consumer",
"chouette",
"chinchin",
"chinaman",
"calderon",
"bullhead",
"brussels",
"brasilia",
"bobby123",
"bellevue",
"bagpipes",
"aurelius",
"altitude",
"aloysius",
"alabama1",
"affinity",
"abcdefg1",
"20102010",
"09876543",
"zxasqw12",
"winnipeg",
"ultraman",
"treefrog",
"tigercat",
"taratara",
"tactical",
"system32",
"swastika",
"skipper1",
"searcher",
"reserved",
"redbeard",
"realtime",
"pyramids",
"provider",
"projects",
"poontang",
"pinecone",
"pericles",
"paradiso",
"parabola",
"overflow",
"mazdarx7",
"marybeth",
"marriott",
"madalena",
"loophole",
"lonsdale",
"lingerie",
"libertad",
"lavalamp",
"joselito",
"joker123",
"jerrylee",
"jamboree",
"interest",
"imissyou",
"hugoboss",
"holahola",
"heythere",
"hehehehe",
"hangover",
"guerrero",
"greatone",
"gianluca",
"gardener",
"gangsta1",
"exorcist",
"dressage",
"dominic1",
"dodgeram",
"cummings",
"christen",
"callahan",
"calcutta",
"burberry",
"betrayal",
"atkinson",
"athletic",
"arachnid",
"amaranth",
"algernon",
"alastair",
"absinthe",
"01020304",
"zoomzoom",
"watchman",
"vanilla1",
"trouble1",
"tortilla",
"squadron",
"smile123",
"skylight",
"ricardo1",
"reliable",
"recorder",
"provence",
"porsche9",
"piedmont",
"patches1",
"overdose",
"nightman",
"mymother",
"monument",
"medicina",
"madonna1",
"longtime",
"lolololo",
"lokiloki",
"laughing",
"kerrigan",
"jeopardy",
"ibelieve",
"houghton",
"horsemen",
"hologram",
"hideaway",
"hawaii50",
"handicap",
"hamsters",
"georgia1",
"freddie1",
"forklift",
"finished",
"dorothea",
"devotion",
"conchita",
"classics",
"chopper1",
"buffalo1",
"bubba123",
"bigballs",
"barnyard",
"baphomet",
"badlands",
"asterisk",
"arcangel",
"20022002",
"19971997",
"whoknows",
"trousers",
"tranquil",
"toriamos",
"temppass",
"teardrop",
"superboy",
"srinivas",
"snowman1",
"shortcut",
"shocking",
"senha123",
"scranton",
"sandoval",
"roseanne",
"red12345",
"prospero",
"products",
"papamama",
"outdoors",
"nemesis1",
"nagasaki",
"mousepad",
"modeling",
"microlab",
"makeitso",
"lalakers",
"kakaroto",
"investor",
"insecure",
"humanoid",
"holiness",
"helpless",
"germaine",
"freefree",
"francais",
"firebolt",
"filipino",
"federica",
"falstaff",
"eleven11",
"dominant",
"diabolic",
"deadbeat",
"crockett",
"crazycat",
"composer",
"coleslaw",
"cascades",
"bretagne",
"breaking",
"bluenose",
"bisexual",
"billions",
"billbill",
"beckham7",
"avengers",
"assembly",
"asasasas",
"allstars",
"alakazam",
"activate",
"Pa55word",
"Computer",
"zerozero",
"vigilant",
"verygood",
"truffles",
"tigerman",
"thankgod",
"telefono",
"summoner",
"suicidal",
"strummer",
"stiletto",
"squeaker",
"sithlord",
"showcase",
"serenade",
"rotation",
"rockhard",
"quintana",
"pacifica",
"omsairam",
"newhouse",
"nacional",
"muenchen",
"morrigan",
"michael2",
"memememe",
"maximize",
"marino13",
"marciano",
"loveable",
"lakeview",
"kenneth1",
"ilikepie",
"historia",
"hiawatha",
"freeport",
"flathead",
"faulkner",
"endymion",
"emirates",
"dreamers",
"dragon69",
"district",
"dietrich",
"clemence",
"claudia1",
"cellular",
"catherin",
"carmella",
"burgundy",
"brother1",
"blooming",
"bigboobs",
"beachbum",
"barbara1",
"backyard",
"backward",
"babybear",
"argonaut",
"appleton",
"aguilera",
"Nicholas",
"Michael1",
"1qazzaq1",
"13243546",
"12qw34er",
"123456ab",
"zaragoza",
"woodcock",
"wisteria",
"westlake",
"victoire",
"trapdoor",
"tigereye",
"thetruth",
"testicle",
"student1",
"sprinkle",
"silencer",
"scottish",
"richelle",
"religion",
"queenbee",
"physical",
"pedersen",
"paperboy",
"nikolaus",
"murderer",
"montague",
"milagros",
"mercutio",
"mercurio",
"mcknight",
"maxpayne",
"manager1",
"mamacita",
"lucretia",
"lol12345",
"laura123",
"kusanagi",
"katmandu",
"julianne",
"joseluis",
"jiujitsu",
"jeanpaul",
"infrared",
"humanity",
"honeypot",
"honeybun",
"herkules",
"hawkeyes",
"gregory1",
"geometry",
"friedman",
"freiheit",
"firework",
"elbereth",
"dragon99",
"dollface",
"devilish",
"democrat",
"darkmoon",
"crackpot",
"costanza",
"consuelo",
"clarisse",
"citibank",
"cingular",
"chrystal",
"channing",
"carvalho",
"brownie1",
"bluebear",
"billyjoe",
"benedikt",
"beaufort",
"batman12",
"barnabas",
"baracuda",
"armitage",
"alcapone",
"adrianne",
"a1a2a3a4",
"Internet",
"Football",
"yourself",
"yorktown",
"yeahyeah",
"valdemar",
"unlocked",
"twinkles",
"trujillo",
"torrents",
"tonyhawk",
"tanzania",
"takedown",
"takamine",
"stitches",
"standing",
"srilanka",
"sparhawk",
"slowpoke",
"shoelace",
"service1",
"senorita",
"seashore",
"roulette",
"rocky123",
"radiator",
"problems",
"platform",
"parallax",
"nepenthe",
"moonmoon",
"lovehate",
"komputer",
"intrigue",
"interact",
"galloway",
"fullback",
"fuckhead",
"fairview",
"divorced",
"disabled",
"defiance",
"deeznutz",
"daniel01",
"cookies1",
"cheating",
"boarding",
"baseline",
"baldrick",
"apollo11",
"aluminum",
"19931993",
"19791979",
"woodwind",
"woodbury",
"watchdog",
"vikings1",
"tribunal",
"toreador",
"thinkpad",
"thebeach",
"terrific",
"teaching",
"stringer",
"souvenir",
"sombrero",
"sk8board",
"shuriken",
"shotokan",
"shinichi",
"scooters",
"regiment",
"rainfall",
"qwerty78",
"pistache",
"pianoman",
"overseas",
"orthodox",
"monorail",
"minemine",
"milhouse",
"mermaids",
"madrigal",
"london22",
"krakatoa",
"junction",
"intranet",
"humility",
"harmless",
"grace123",
"giuliana",
"gauntlet",
"fugitive",
"flatland",
"feelings",
"fabregas",
"emanuele",
"election",
"dumpster",
"douglas1",
"cruzeiro",
"cracking",
"control1",
"cheaters",
"centrino",
"captain1",
"canberra",
"botswana",
"atreides",
"asuncion",
"astroboy",
"aqualung",
"amnesiac",
"adorable",
"3edc4rfv",
"1z2x3c4v",
"19921992",
"14141414",
"12211221",
"yankees2",
"worldcup",
"vittorio",
"theworld",
"thebeast",
"thaddeus",
"telemark",
"sylvania",
"surveyor",
"suitcase",
"stroller",
"stripped",
"stallone",
"smoke420",
"septembe",
"sandberg",
"rousseau",
"revenant",
"pepsi123",
"pembroke",
"parkside",
"outbreak",
"obsolete",
"nutshell",
"nounours",
"nonenone",
"momentum",
"michele1",
"maldives",
"magdalen",
"lockhart",
"krokodil",
"humboldt",
"homebase",
"headshot",
"headless",
"hazelnut",
"gremlins",
"frankie1",
"frank123",
"fireman1",
"external",
"entering",
"dulcinea",
"dropkick",
"draconis",
"dont4get",
"domestic",
"darkwing",
"corporal",
"cocorico",
"chimaera",
"cheyanne",
"breakers",
"bluesman",
"bethesda",
"basketba",
"andyandy",
"allison1",
"Garfield",
"Abcd1234",
"yoyoyoyo",
"yeahbaby",
"wetpussy",
"variable",
"unicorn1",
"trillium",
"torrance",
"tikitiki",
"thumper1",
"thesaint",
"theforce",
"teiubesc",
"sweet123",
"succubus",
"stockman",
"steve123",
"speeding",
"sokrates",
"showboat",
"sequence",
"qwerty99",
"postcard",
"polkadot",
"orlando1",
"nicolas1",
"nicknick",
"naughty1",
"marielle",
"maneater",
"lionlion",
"leapfrog",
"kirkwood",
"kilkenny",
"jordan12",
"intercom",
"informix",
"hounddog",
"homicide",
"herschel",
"hatteras",
"harakiri",
"halfmoon",
"fivestar",
"firewood",
"executor",
"elcamino",
"egyptian",
"eclipse1",
"duckling",
"drumming",
"drifting",
"daisydog",
"coolgirl",
"contrast",
"choclate",
"chilling",
"channels",
"catapult",
"careless",
"californ",
"brendan1",
"beverley",
"atalanta",
"ashley12",
"arizona1",
"antihero",
"andrew12",
"allright",
"ab123456",
"43214321",
"18436572",
"windows7",
"wellcome",
"waldemar",
"valerian",
"tristan1",
"tornado1",
"thunders",
"tennyson",
"tarragon",
"tapestry",
"tajmahal",
"sunny123",
"struggle",
"starling",
"sobriety",
"snowfall",
"skyline1",
"shirley1",
"shalimar",
"settings",
"schnecke",
"satriani",
"sasha123",
"sailfish",
"roserose",
"qwerty22",
"prashant",
"powerman",
"powerade",
"plastics",
"pinkpink",
"parallel",
"papercut",
"p4ssword",
"navyseal",
"monopoli",
"mnemonic",
"millenia",
"membrane",
"manitoba",
"lineage2",
"leopards",
"karoline",
"johnpaul",
"interior",
"homepage",
"greeting",
"golfgolf",
"glassman",
"friction",
"filomena",
"ethereal",
"emotions",
"dudedude",
"douglass",
"dominika",
"demetrio",
"demented",
"decision",
"cuthbert",
"compound",
"comatose",
"civilwar",
"castello",
"cachorro",
"bulletin",
"brandnew",
"bluegill",
"baywatch",
"bastardo",
"bagheera",
"annalisa",
"allstate",
"alberto1",
"Samantha",
"78945612",
"01010101",
"yellow12",
"wildbill",
"whittier",
"vittoria",
"virgilio",
"trusting",
"troubles",
"tonytony",
"thebest1",
"terriers",
"template",
"telefoon",
"talented",
"supermen",
"starting",
"sixpence",
"sidewalk",
"shoshana",
"rainbow7",
"rafferty",
"qwerty77",
"qwerty00",
"pheasant",
"pentium3",
"patrizia",
"overlook",
"overhead",
"okokokok",
"nwo4life",
"novembre",
"newlife1",
"newdelhi",
"myspace1",
"myfriend",
"munchies",
"moneybag",
"molecule",
"mercury1",
"melville",
"mcintyre",
"mattress",
"maritime",
"mariachi",
"loveyou2",
"lovesong",
"lolalola",
"lindsey1",
"lifeboat",
"katie123",
"kasandra",
"jupiter1",
"julia123",
"india123",
"henry123",
"henrique",
"hardball",
"handbook",
"hacienda",
"grenoble",
"giuliano",
"freehand",
"fragment",
"foreskin",
"ensemble",
"eclectic",
"dogfight",
"dodgers1",
"diogenes",
"dillweed",
"demon666",
"daybreak",
"dagobert",
"culinary",
"crossing",
"controls",
"cobblers",
"charissa",
"buster12",
"bungalow",
"brianna1",
"bella123",
"ballroom",
"andre123",
"analysis",
"amber123",
"aa123456",
"2wsx3edc",
"12131213",
"wertwert",
"vivienne",
"tuppence",
"trafford",
"teddy123",
"streamer",
"star1234",
"sparrows",
"solomon1",
"sideshow",
"sherbert",
"sebastia",
"scribble",
"sarasota",
"sarasara",
"sarah123",
"sanguine",
"sandy123",
"robert12",
"redhorse",
"rational",
"radioman",
"qwerty01",
"poophead",
"phantoms",
"paperino",
"organize",
"optiplex",
"october1",
"neverdie",
"monsieur",
"monkfish",
"master01",
"marymary",
"lucas123",
"logistic",
"lemmings",
"langston",
"killer11",
"jack1234",
"ireland1",
"house123",
"hihihihi",
"hellhole",
"hardwood",
"funhouse",
"fiorella",
"farewell",
"fantasma",
"failsafe",
"explicit",
"esposito",
"duckduck",
"drilling",
"dragon10",
"dickweed",
"crunchie",
"crawfish",
"chessman",
"chanelle",
"chamonix",
"candy123",
"brainiac",
"birdland",
"binladen",
"billings",
"bareback",
"bacteria",
"asdfqwer",
"asd12345",
"arpeggio",
"anthony2",
"animator",
"amazonas",
"alpacino",
"adelaida",
"adamadam",
"aaron123",
"Einstein",
"90909090",
"1234zxcv",
"yamamoto",
"wormhole",
"whiteman",
"westgate",
"watchmen",
"vergeten",
"veracruz",
"vanquish",
"uuuuuuuu",
"trucking",
"trooper1",
"timelord",
"strangle",
"stoneman",
"starless",
"spagetti",
"sorensen",
"somethin",
"snowhite",
"slovakia",
"skydiver",
"silicone",
"silencio",
"selector",
"scramble",
"scott123",
"salinger",
"reminder",
"redheads",
"phaedrus",
"paulchen",
"passion1",
"paraguay",
"panda123",
"palacios",
"osbourne",
"onepiece",
"mutation",
"murakami",
"mercator",
"mario123",
"lynnette",
"lookatme",
"linda123",
"lightnin",
"lifeless",
"leopoldo",
"kristin1",
"knitting",
"katrina1",
"hershey1",
"gridlock",
"gigantic",
"fred1234",
"flatline",
"firehawk",
"fellatio",
"eruption",
"dragons1",
"dragon88",
"delorean",
"decipher",
"darkblue",
"creatine",
"counting",
"coolidge",
"cookie12",
"converge",
"clubbing",
"cbr600rr",
"carnegie",
"calabria",
"buttfuck",
"broncos1",
"blueball",
"beautifu",
"barnacle",
"babygurl",
"asturias",
"armchair",
"archives",
"aperture",
"amandine",
"22446688",
"20032003",
"19641964",
"12141214",
"01230123",
"yourname",
"warszawa",
"therock1",
"testuser",
"temp1234",
"swordfis",
"superdog",
"sunflowe",
"soccer22",
"slovenia",
"sinfonia",
"scimitar",
"rosebush",
"redriver",
"redeemed",
"ramstein",
"qweasdzx",
"plumbing",
"pickwick",
"parsifal",
"overcome",
"ninjutsu",
"newport1",
"newcomer",
"monkey01",
"minority",
"mariette",
"loveland",
"lagrange",
"kaitlynn",
"john1234",
"invictus",
"inventor",
"inspired",
"hurrican",
"honey123",
"holbrook",
"heracles",
"hathaway",
"governor",
"goodrich",
"gizmo123",
"friday13",
"fortytwo",
"foreplay",
"fishhook",
"fishfish",
"fillmore",
"espinoza",
"emerald1",
"edgewood",
"duisburg",
"drummers",
"dowjones",
"cameroon",
"buddyboy",
"bracelet",
"bogeyman",
"bluerose",
"birdcage",
"billy123",
"beepbeep",
"asdfgh12",
"antonina",
"anabolic",
"allister",
"albacore",
"airedale",
"activity",
"Patricia",
"99887766",
"20202020",
"19701970",
"yardbird",
"xcountry",
"wildrose",
"watanabe",
"wareagle",
"validate",
"tripping",
"treetree",
"timbuktu",
"summer00",
"stuntman",
"steelman",
"spartan1",
"snowshoe",
"smuggler",
"slowhand",
"shadow01",
"schuster",
"satelite",
"rightnow",
"r4e3w2q1",
"quagmire",
"porridge",
"peerless",
"paganini",
"optional",
"nowayout",
"newstart",
"neworder",
"monkey13",
"mission1",
"mcmillan",
"lucky777",
"lombardo",
"lindberg",
"larkspur",
"lambchop",
"lalaland",
"kirakira",
"joshua12",
"january1",
"infinito",
"identify",
"hellgate",
"heatwave",
"grounded",
"greenish",
"gorillaz",
"gerhardt",
"generous",
"gauthier",
"frontera",
"freezing",
"fracture",
"fastlane",
"drafting",
"donnelly",
"dolomite",
"damocles",
"critters",
"crickets",
"crabtree",
"cortland",
"comrades",
"clothing",
"checking",
"charmed1",
"cathleen",
"carter15",
"carleton",
"blueline",
"bigblack",
"bastard1",
"backspin",
"babababa",
"audition",
"argentum",
"antonius",
"antiques",
"abigail1",
"14531453",
"woodlawn",
"windward",
"warranty",
"visitors",
"trespass",
"trashcan",
"topnotch",
"tigger12",
"summer05",
"summer01",
"sturgeon",
"strikers",
"skipjack",
"shipyard",
"shekinah",
"scouting",
"sanpedro",
"sandrock",
"rootroot",
"ronaldo9",
"reynaldo",
"relative",
"radagast",
"qwertzui",
"presidio",
"presence",
"prentice",
"playback",
"philippa",
"peterman",
"peregrin",
"peaceman",
"papabear",
"organist",
"octavian",
"nascar24",
"monteiro",
"monkeys1",
"metaphor",
"manifold",
"makelove",
"lysander",
"lobsters",
"julie123",
"johngalt",
"jamaica1",
"jalapeno",
"jacobsen",
"isengard",
"hutchins",
"horizons",
"hawkwind",
"happyboy",
"gutentag",
"gracious",
"glenwood",
"frogfrog",
"fraction",
"folklore",
"fantasy1",
"express1",
"exposure",
"everton1",
"employee",
"economic",
"ducksoup",
"diskette",
"delacruz",
"creepers",
"clements",
"cheerful",
"catering",
"capucine",
"capacity",
"bridgett",
"boyscout",
"bingo123",
"belgrade",
"beginner",
"bavarian",
"backfire",
"astaroth",
"arsehole",
"annelise",
"andrew01",
"anabelle",
"albright",
"airlines",
"adelante",
"account1",
"Maverick",
"85208520",
"14121412",
"yahoo123",
"wretched",
"winthrop",
"westwind",
"weinberg",
"trashman",
"toronto1",
"thomas01",
"thibault",
"syndrome",
"swinging",
"sweetest",
"sunburst",
"sperling",
"spectral",
"soldier1",
"silmaril",
"shoulder",
"shahrukh",
"settlers",
"scotsman",
"scofield",
"schumann",
"rockrock",
"rockland",
"qwerty69",
"promises",
"priscila",
"priority",
"playoffs",
"pebbles1",
"overseer",
"opposite",
"octavius",
"nikenike",
"nehemiah",
"mystery1",
"morticia",
"monkey11",
"misty123",
"milenium",
"michael3",
"lincoln1",
"lilwayne",
"lausanne",
"kokokoko",
"kilowatt",
"jacob123",
"interval",
"ignorant",
"huntsman",
"homesick",
"highbury",
"hellbent",
"guerilla",
"graywolf",
"grandson",
"gargamel",
"gameplay",
"firefly1",
"fighter1",
"fielding",
"familiar",
"falconer",
"ezequiel",
"dynamics",
"demetria",
"darkroom",
"curtains",
"currency",
"crocodil",
"crawling",
"christy1",
"chivalry",
"charlie7",
"catriona",
"carolann",
"cantona7",
"canfield",
"buttocks",
"brinkley",
"bordello",
"blissful",
"blackbox",
"billiard",
"bigbooty",
"bastille",
"as123456",
"artofwar",
"annalena",
"animated",
"alvarado",
"alicante",
"alex2000",
"accurate",
"17171717",
"123456as",
"00112233",
"00001111"
};